module heichips25_top_sorter (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire \s0.data_new_delayed[0] ;
 wire \s0.data_new_delayed[1] ;
 wire \s0.data_new_delayed[2] ;
 wire \s0.data_new_delayed[3] ;
 wire \s0.data_new_delayed[4] ;
 wire \s0.data_new_delayed[5] ;
 wire \s0.data_new_delayed[6] ;
 wire \s0.data_new_delayed[7] ;
 wire \s0.data_out[0][0] ;
 wire \s0.data_out[0][1] ;
 wire \s0.data_out[0][2] ;
 wire \s0.data_out[0][3] ;
 wire \s0.data_out[0][4] ;
 wire \s0.data_out[0][5] ;
 wire \s0.data_out[0][6] ;
 wire \s0.data_out[0][7] ;
 wire \s0.data_out[10][0] ;
 wire \s0.data_out[10][1] ;
 wire \s0.data_out[10][2] ;
 wire \s0.data_out[10][3] ;
 wire \s0.data_out[10][4] ;
 wire \s0.data_out[10][5] ;
 wire \s0.data_out[10][6] ;
 wire \s0.data_out[10][7] ;
 wire \s0.data_out[11][0] ;
 wire \s0.data_out[11][1] ;
 wire \s0.data_out[11][2] ;
 wire \s0.data_out[11][3] ;
 wire \s0.data_out[11][4] ;
 wire \s0.data_out[11][5] ;
 wire \s0.data_out[11][6] ;
 wire \s0.data_out[11][7] ;
 wire \s0.data_out[12][0] ;
 wire \s0.data_out[12][1] ;
 wire \s0.data_out[12][2] ;
 wire \s0.data_out[12][3] ;
 wire \s0.data_out[12][4] ;
 wire \s0.data_out[12][5] ;
 wire \s0.data_out[12][6] ;
 wire \s0.data_out[12][7] ;
 wire \s0.data_out[13][0] ;
 wire \s0.data_out[13][1] ;
 wire \s0.data_out[13][2] ;
 wire \s0.data_out[13][3] ;
 wire \s0.data_out[13][4] ;
 wire \s0.data_out[13][5] ;
 wire \s0.data_out[13][6] ;
 wire \s0.data_out[13][7] ;
 wire \s0.data_out[14][0] ;
 wire \s0.data_out[14][1] ;
 wire \s0.data_out[14][2] ;
 wire \s0.data_out[14][3] ;
 wire \s0.data_out[14][4] ;
 wire \s0.data_out[14][5] ;
 wire \s0.data_out[14][6] ;
 wire \s0.data_out[14][7] ;
 wire \s0.data_out[15][0] ;
 wire \s0.data_out[15][1] ;
 wire \s0.data_out[15][2] ;
 wire \s0.data_out[15][3] ;
 wire \s0.data_out[15][4] ;
 wire \s0.data_out[15][5] ;
 wire \s0.data_out[15][6] ;
 wire \s0.data_out[15][7] ;
 wire \s0.data_out[16][0] ;
 wire \s0.data_out[16][1] ;
 wire \s0.data_out[16][2] ;
 wire \s0.data_out[16][3] ;
 wire \s0.data_out[16][4] ;
 wire \s0.data_out[16][5] ;
 wire \s0.data_out[16][6] ;
 wire \s0.data_out[16][7] ;
 wire \s0.data_out[17][0] ;
 wire \s0.data_out[17][1] ;
 wire \s0.data_out[17][2] ;
 wire \s0.data_out[17][3] ;
 wire \s0.data_out[17][4] ;
 wire \s0.data_out[17][5] ;
 wire \s0.data_out[17][6] ;
 wire \s0.data_out[17][7] ;
 wire \s0.data_out[18][0] ;
 wire \s0.data_out[18][1] ;
 wire \s0.data_out[18][2] ;
 wire \s0.data_out[18][3] ;
 wire \s0.data_out[18][4] ;
 wire \s0.data_out[18][5] ;
 wire \s0.data_out[18][6] ;
 wire \s0.data_out[18][7] ;
 wire \s0.data_out[19][0] ;
 wire \s0.data_out[19][1] ;
 wire \s0.data_out[19][2] ;
 wire \s0.data_out[19][3] ;
 wire \s0.data_out[19][4] ;
 wire \s0.data_out[19][5] ;
 wire \s0.data_out[19][6] ;
 wire \s0.data_out[19][7] ;
 wire \s0.data_out[1][0] ;
 wire \s0.data_out[1][1] ;
 wire \s0.data_out[1][2] ;
 wire \s0.data_out[1][3] ;
 wire \s0.data_out[1][4] ;
 wire \s0.data_out[1][5] ;
 wire \s0.data_out[1][6] ;
 wire \s0.data_out[1][7] ;
 wire \s0.data_out[20][0] ;
 wire \s0.data_out[20][1] ;
 wire \s0.data_out[20][2] ;
 wire \s0.data_out[20][3] ;
 wire \s0.data_out[20][4] ;
 wire \s0.data_out[20][5] ;
 wire \s0.data_out[20][6] ;
 wire \s0.data_out[20][7] ;
 wire \s0.data_out[21][0] ;
 wire \s0.data_out[21][1] ;
 wire \s0.data_out[21][2] ;
 wire \s0.data_out[21][3] ;
 wire \s0.data_out[21][4] ;
 wire \s0.data_out[21][5] ;
 wire \s0.data_out[21][6] ;
 wire \s0.data_out[21][7] ;
 wire \s0.data_out[2][0] ;
 wire \s0.data_out[2][1] ;
 wire \s0.data_out[2][2] ;
 wire \s0.data_out[2][3] ;
 wire \s0.data_out[2][4] ;
 wire \s0.data_out[2][5] ;
 wire \s0.data_out[2][6] ;
 wire \s0.data_out[2][7] ;
 wire \s0.data_out[3][0] ;
 wire \s0.data_out[3][1] ;
 wire \s0.data_out[3][2] ;
 wire \s0.data_out[3][3] ;
 wire \s0.data_out[3][4] ;
 wire \s0.data_out[3][5] ;
 wire \s0.data_out[3][6] ;
 wire \s0.data_out[3][7] ;
 wire \s0.data_out[4][0] ;
 wire \s0.data_out[4][1] ;
 wire \s0.data_out[4][2] ;
 wire \s0.data_out[4][3] ;
 wire \s0.data_out[4][4] ;
 wire \s0.data_out[4][5] ;
 wire \s0.data_out[4][6] ;
 wire \s0.data_out[4][7] ;
 wire \s0.data_out[5][0] ;
 wire \s0.data_out[5][1] ;
 wire \s0.data_out[5][2] ;
 wire \s0.data_out[5][3] ;
 wire \s0.data_out[5][4] ;
 wire \s0.data_out[5][5] ;
 wire \s0.data_out[5][6] ;
 wire \s0.data_out[5][7] ;
 wire \s0.data_out[6][0] ;
 wire \s0.data_out[6][1] ;
 wire \s0.data_out[6][2] ;
 wire \s0.data_out[6][3] ;
 wire \s0.data_out[6][4] ;
 wire \s0.data_out[6][5] ;
 wire \s0.data_out[6][6] ;
 wire \s0.data_out[6][7] ;
 wire \s0.data_out[7][0] ;
 wire \s0.data_out[7][1] ;
 wire \s0.data_out[7][2] ;
 wire \s0.data_out[7][3] ;
 wire \s0.data_out[7][4] ;
 wire \s0.data_out[7][5] ;
 wire \s0.data_out[7][6] ;
 wire \s0.data_out[7][7] ;
 wire \s0.data_out[8][0] ;
 wire \s0.data_out[8][1] ;
 wire \s0.data_out[8][2] ;
 wire \s0.data_out[8][3] ;
 wire \s0.data_out[8][4] ;
 wire \s0.data_out[8][5] ;
 wire \s0.data_out[8][6] ;
 wire \s0.data_out[8][7] ;
 wire \s0.data_out[9][0] ;
 wire \s0.data_out[9][1] ;
 wire \s0.data_out[9][2] ;
 wire \s0.data_out[9][3] ;
 wire \s0.data_out[9][4] ;
 wire \s0.data_out[9][5] ;
 wire \s0.data_out[9][6] ;
 wire \s0.data_out[9][7] ;
 wire \s0.genblk1[10].modules.bubble ;
 wire \s0.genblk1[11].modules.bubble ;
 wire \s0.genblk1[12].modules.bubble ;
 wire \s0.genblk1[13].modules.bubble ;
 wire \s0.genblk1[14].modules.bubble ;
 wire \s0.genblk1[15].modules.bubble ;
 wire \s0.genblk1[16].modules.bubble ;
 wire \s0.genblk1[17].modules.bubble ;
 wire \s0.genblk1[18].modules.bubble ;
 wire \s0.genblk1[19].modules.bubble ;
 wire \s0.genblk1[1].modules.bubble ;
 wire \s0.genblk1[20].modules.bubble ;
 wire \s0.genblk1[21].modules.bubble ;
 wire \s0.genblk1[2].modules.bubble ;
 wire \s0.genblk1[3].modules.bubble ;
 wire \s0.genblk1[4].modules.bubble ;
 wire \s0.genblk1[5].modules.bubble ;
 wire \s0.genblk1[6].modules.bubble ;
 wire \s0.genblk1[7].modules.bubble ;
 wire \s0.genblk1[8].modules.bubble ;
 wire \s0.genblk1[9].modules.bubble ;
 wire \s0.module0.bubble ;
 wire net11;
 wire net12;
 wire net296;
 wire net13;
 wire net14;
 wire clknet_leaf_0_clk;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net1;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net10;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire [0:0] \s0.shift_out[0] ;
 wire [0:0] \s0.shift_out[10] ;
 wire [0:0] \s0.shift_out[11] ;
 wire [0:0] \s0.shift_out[12] ;
 wire [0:0] \s0.shift_out[13] ;
 wire [0:0] \s0.shift_out[14] ;
 wire [0:0] \s0.shift_out[15] ;
 wire [0:0] \s0.shift_out[16] ;
 wire [0:0] \s0.shift_out[17] ;
 wire [0:0] \s0.shift_out[18] ;
 wire [0:0] \s0.shift_out[19] ;
 wire [0:0] \s0.shift_out[1] ;
 wire [0:0] \s0.shift_out[20] ;
 wire [0:0] \s0.shift_out[21] ;
 wire [0:0] \s0.shift_out[2] ;
 wire [0:0] \s0.shift_out[3] ;
 wire [0:0] \s0.shift_out[4] ;
 wire [0:0] \s0.shift_out[5] ;
 wire [0:0] \s0.shift_out[6] ;
 wire [0:0] \s0.shift_out[7] ;
 wire [0:0] \s0.shift_out[8] ;
 wire [0:0] \s0.shift_out[9] ;
 wire [0:0] \s0.valid_out[0] ;
 wire [0:0] \s0.valid_out[10] ;
 wire [0:0] \s0.valid_out[11] ;
 wire [0:0] \s0.valid_out[12] ;
 wire [0:0] \s0.valid_out[13] ;
 wire [0:0] \s0.valid_out[14] ;
 wire [0:0] \s0.valid_out[15] ;
 wire [0:0] \s0.valid_out[16] ;
 wire [0:0] \s0.valid_out[17] ;
 wire [0:0] \s0.valid_out[18] ;
 wire [0:0] \s0.valid_out[19] ;
 wire [0:0] \s0.valid_out[1] ;
 wire [0:0] \s0.valid_out[20] ;
 wire [0:0] \s0.valid_out[21] ;
 wire [0:0] \s0.valid_out[2] ;
 wire [0:0] \s0.valid_out[3] ;
 wire [0:0] \s0.valid_out[4] ;
 wire [0:0] \s0.valid_out[5] ;
 wire [0:0] \s0.valid_out[6] ;
 wire [0:0] \s0.valid_out[7] ;
 wire [0:0] \s0.valid_out[8] ;
 wire [0:0] \s0.valid_out[9] ;
 wire [0:0] \s0.was_valid_out[0] ;
 wire [0:0] \s0.was_valid_out[10] ;
 wire [0:0] \s0.was_valid_out[11] ;
 wire [0:0] \s0.was_valid_out[12] ;
 wire [0:0] \s0.was_valid_out[13] ;
 wire [0:0] \s0.was_valid_out[14] ;
 wire [0:0] \s0.was_valid_out[15] ;
 wire [0:0] \s0.was_valid_out[16] ;
 wire [0:0] \s0.was_valid_out[17] ;
 wire [0:0] \s0.was_valid_out[18] ;
 wire [0:0] \s0.was_valid_out[19] ;
 wire [0:0] \s0.was_valid_out[1] ;
 wire [0:0] \s0.was_valid_out[20] ;
 wire [0:0] \s0.was_valid_out[21] ;
 wire [0:0] \s0.was_valid_out[2] ;
 wire [0:0] \s0.was_valid_out[3] ;
 wire [0:0] \s0.was_valid_out[4] ;
 wire [0:0] \s0.was_valid_out[5] ;
 wire [0:0] \s0.was_valid_out[6] ;
 wire [0:0] \s0.was_valid_out[7] ;
 wire [0:0] \s0.was_valid_out[8] ;
 wire [0:0] \s0.was_valid_out[9] ;

 sg13g2_nand2_1 _3107_ (.Y(_1564_),
    .A(net1020),
    .B(net411));
 sg13g2_mux2_1 _3108_ (.A0(\s0.data_out[8][4] ),
    .A1(\s0.data_out[7][4] ),
    .S(net1021),
    .X(_1565_));
 sg13g2_a21oi_1 _3109_ (.A1(net1016),
    .A2(_1565_),
    .Y(_1566_),
    .B1(_1508_));
 sg13g2_nand2b_1 _3110_ (.Y(_1567_),
    .B(net1025),
    .A_N(_1566_));
 sg13g2_nand3_1 _3111_ (.B(_1506_),
    .C(_1567_),
    .A(net1256),
    .Y(_1568_));
 sg13g2_nand2_1 _3112_ (.Y(_1569_),
    .A(net1020),
    .B(net589));
 sg13g2_mux2_1 _3113_ (.A0(\s0.data_out[8][5] ),
    .A1(\s0.data_out[7][5] ),
    .S(net1021),
    .X(_1570_));
 sg13g2_a21o_1 _3114_ (.A2(_1570_),
    .A1(net1016),
    .B1(_1514_),
    .X(_1571_));
 sg13g2_a21oi_1 _3115_ (.A1(net1026),
    .A2(_1571_),
    .Y(_1572_),
    .B1(_1513_));
 sg13g2_nand2_1 _3116_ (.Y(_1573_),
    .A(net1252),
    .B(_1572_));
 sg13g2_a21o_1 _3117_ (.A2(_1567_),
    .A1(_1506_),
    .B1(net1256),
    .X(_1574_));
 sg13g2_nor2_1 _3118_ (.A(net1252),
    .B(_1572_),
    .Y(_1575_));
 sg13g2_o21ai_1 _3119_ (.B1(_1573_),
    .Y(_1576_),
    .A1(net1266),
    .A2(_1549_));
 sg13g2_nor3_1 _3120_ (.A(_1563_),
    .B(_1575_),
    .C(_1576_),
    .Y(_1577_));
 sg13g2_nand4_1 _3121_ (.B(_1568_),
    .C(_1574_),
    .A(_1551_),
    .Y(_1578_),
    .D(_1577_));
 sg13g2_o21ai_1 _3122_ (.B1(_1573_),
    .Y(_1579_),
    .A1(_1568_),
    .A2(_1575_));
 sg13g2_nor2b_1 _3123_ (.A(_1563_),
    .B_N(_1579_),
    .Y(_1580_));
 sg13g2_nor2b_1 _3124_ (.A(_1560_),
    .B_N(_1562_),
    .Y(_1581_));
 sg13g2_nor3_1 _3125_ (.A(_1471_),
    .B(_1580_),
    .C(_1581_),
    .Y(_1582_));
 sg13g2_or2_1 _3126_ (.X(_1583_),
    .B(net1209),
    .A(net307));
 sg13g2_a21oi_1 _3127_ (.A1(_1578_),
    .A2(_1582_),
    .Y(_0174_),
    .B1(_1583_));
 sg13g2_and2_1 _3128_ (.A(net1326),
    .B(net313),
    .X(_0175_));
 sg13g2_o21ai_1 _3129_ (.B1(net1015),
    .Y(_1584_),
    .A1(net1228),
    .A2(net1005));
 sg13g2_nor2b_1 _3130_ (.A(net1228),
    .B_N(net1010),
    .Y(_1585_));
 sg13g2_nor2_1 _3131_ (.A(_1584_),
    .B(_1585_),
    .Y(_1586_));
 sg13g2_o21ai_1 _3132_ (.B1(_1586_),
    .Y(_1587_),
    .A1(\s0.was_valid_out[6] [0]),
    .A2(net1010));
 sg13g2_nor2_1 _3133_ (.A(net1005),
    .B(_1584_),
    .Y(_1588_));
 sg13g2_o21ai_1 _3134_ (.B1(_2468_),
    .Y(_1589_),
    .A1(\s0.was_valid_out[6] [0]),
    .A2(net1020));
 sg13g2_nand2_1 _3135_ (.Y(_1590_),
    .A(_1587_),
    .B(_1589_));
 sg13g2_a21oi_1 _3136_ (.A1(net1222),
    .A2(net1020),
    .Y(_1591_),
    .B1(net1015));
 sg13g2_nor2_1 _3137_ (.A(_1586_),
    .B(_1591_),
    .Y(_1592_));
 sg13g2_o21ai_1 _3138_ (.B1(net1329),
    .Y(_1593_),
    .A1(_1588_),
    .A2(_1590_));
 sg13g2_a21oi_1 _3139_ (.A1(_2444_),
    .A2(_1592_),
    .Y(_0176_),
    .B1(_1593_));
 sg13g2_nor3_1 _3140_ (.A(net1220),
    .B(_1586_),
    .C(_1591_),
    .Y(_0177_));
 sg13g2_mux2_1 _3141_ (.A0(\s0.data_out[6][0] ),
    .A1(\s0.data_out[7][0] ),
    .S(net1019),
    .X(_1594_));
 sg13g2_nand2_1 _3142_ (.Y(_1595_),
    .A(net917),
    .B(_1594_));
 sg13g2_and2_1 _3143_ (.A(net1001),
    .B(\s0.data_out[6][0] ),
    .X(_1596_));
 sg13g2_nor2b_1 _3144_ (.A(net1001),
    .B_N(net1074),
    .Y(_1597_));
 sg13g2_o21ai_1 _3145_ (.B1(net1012),
    .Y(_1598_),
    .A1(_1596_),
    .A2(_1597_));
 sg13g2_nand3_1 _3146_ (.B(_1595_),
    .C(_1598_),
    .A(net1327),
    .Y(_1599_));
 sg13g2_o21ai_1 _3147_ (.B1(_1599_),
    .Y(_1600_),
    .A1(net1327),
    .A2(net391));
 sg13g2_inv_1 _3148_ (.Y(_0178_),
    .A(_1600_));
 sg13g2_mux2_1 _3149_ (.A0(\s0.data_out[6][1] ),
    .A1(\s0.data_out[7][1] ),
    .S(net1019),
    .X(_1601_));
 sg13g2_nand2_1 _3150_ (.Y(_1602_),
    .A(net917),
    .B(_1601_));
 sg13g2_and2_1 _3151_ (.A(net1001),
    .B(\s0.data_out[6][1] ),
    .X(_1603_));
 sg13g2_nor2b_1 _3152_ (.A(net1002),
    .B_N(net1071),
    .Y(_1604_));
 sg13g2_o21ai_1 _3153_ (.B1(net1012),
    .Y(_1605_),
    .A1(_1603_),
    .A2(_1604_));
 sg13g2_nand3_1 _3154_ (.B(_1602_),
    .C(_1605_),
    .A(net1327),
    .Y(_1606_));
 sg13g2_o21ai_1 _3155_ (.B1(_1606_),
    .Y(_1607_),
    .A1(net1327),
    .A2(net419));
 sg13g2_inv_1 _3156_ (.Y(_0179_),
    .A(_1607_));
 sg13g2_mux2_1 _3157_ (.A0(\s0.data_out[6][2] ),
    .A1(\s0.data_out[7][2] ),
    .S(net1019),
    .X(_1608_));
 sg13g2_nand2_1 _3158_ (.Y(_1609_),
    .A(net917),
    .B(_1608_));
 sg13g2_and2_1 _3159_ (.A(net1001),
    .B(\s0.data_out[6][2] ),
    .X(_1610_));
 sg13g2_nor2b_1 _3160_ (.A(net1001),
    .B_N(net1066),
    .Y(_1611_));
 sg13g2_o21ai_1 _3161_ (.B1(net1012),
    .Y(_1612_),
    .A1(_1610_),
    .A2(_1611_));
 sg13g2_nand3_1 _3162_ (.B(_1609_),
    .C(_1612_),
    .A(net1327),
    .Y(_1613_));
 sg13g2_o21ai_1 _3163_ (.B1(_1613_),
    .Y(_1614_),
    .A1(net1324),
    .A2(net467));
 sg13g2_inv_1 _3164_ (.Y(_0180_),
    .A(_1614_));
 sg13g2_nand2b_1 _3165_ (.Y(_1615_),
    .B(net454),
    .A_N(net1019));
 sg13g2_a21oi_1 _3166_ (.A1(_1545_),
    .A2(_1615_),
    .Y(_1616_),
    .B1(net1012));
 sg13g2_nor2b_1 _3167_ (.A(net1002),
    .B_N(net1062),
    .Y(_1617_));
 sg13g2_a21oi_1 _3168_ (.A1(net1002),
    .A2(net454),
    .Y(_1618_),
    .B1(_1617_));
 sg13g2_o21ai_1 _3169_ (.B1(net1327),
    .Y(_1619_),
    .A1(net917),
    .A2(_1618_));
 sg13g2_or2_1 _3170_ (.X(_1620_),
    .B(net503),
    .A(net1327));
 sg13g2_o21ai_1 _3171_ (.B1(_1620_),
    .Y(_1621_),
    .A1(_1616_),
    .A2(_1619_));
 sg13g2_inv_1 _3172_ (.Y(_0181_),
    .A(_1621_));
 sg13g2_nand2b_1 _3173_ (.Y(_1622_),
    .B(net423),
    .A_N(net1019));
 sg13g2_a21oi_1 _3174_ (.A1(_1564_),
    .A2(_1622_),
    .Y(_1623_),
    .B1(net1015));
 sg13g2_nor2b_1 _3175_ (.A(net1005),
    .B_N(net1059),
    .Y(_1624_));
 sg13g2_a21oi_1 _3176_ (.A1(net1005),
    .A2(net423),
    .Y(_1625_),
    .B1(_1624_));
 sg13g2_o21ai_1 _3177_ (.B1(net1329),
    .Y(_1626_),
    .A1(_2468_),
    .A2(_1625_));
 sg13g2_or2_1 _3178_ (.X(_1627_),
    .B(net411),
    .A(net1329));
 sg13g2_o21ai_1 _3179_ (.B1(_1627_),
    .Y(_1628_),
    .A1(_1623_),
    .A2(_1626_));
 sg13g2_inv_1 _3180_ (.Y(_0182_),
    .A(_1628_));
 sg13g2_nand2b_1 _3181_ (.Y(_1629_),
    .B(net539),
    .A_N(net1020));
 sg13g2_a21oi_1 _3182_ (.A1(_1569_),
    .A2(_1629_),
    .Y(_1630_),
    .B1(net1015));
 sg13g2_nor2b_1 _3183_ (.A(net1005),
    .B_N(net1055),
    .Y(_1631_));
 sg13g2_a21oi_1 _3184_ (.A1(net1005),
    .A2(net539),
    .Y(_1632_),
    .B1(_1631_));
 sg13g2_o21ai_1 _3185_ (.B1(net1326),
    .Y(_1633_),
    .A1(_2468_),
    .A2(_1632_));
 sg13g2_or2_1 _3186_ (.X(_1634_),
    .B(net589),
    .A(net1329));
 sg13g2_o21ai_1 _3187_ (.B1(_1634_),
    .Y(_1635_),
    .A1(_1630_),
    .A2(_1633_));
 sg13g2_inv_1 _3188_ (.Y(_0183_),
    .A(_1635_));
 sg13g2_nand2b_1 _3189_ (.Y(_1636_),
    .B(\s0.data_out[6][6] ),
    .A_N(net1020));
 sg13g2_a21oi_1 _3190_ (.A1(_1556_),
    .A2(_1636_),
    .Y(_1637_),
    .B1(net1015));
 sg13g2_nor2b_1 _3191_ (.A(net1006),
    .B_N(net1051),
    .Y(_1638_));
 sg13g2_a21oi_1 _3192_ (.A1(net1006),
    .A2(\s0.data_out[6][6] ),
    .Y(_1639_),
    .B1(_1638_));
 sg13g2_o21ai_1 _3193_ (.B1(net1326),
    .Y(_1640_),
    .A1(net917),
    .A2(_1639_));
 sg13g2_or2_1 _3194_ (.X(_1641_),
    .B(net544),
    .A(net1329));
 sg13g2_o21ai_1 _3195_ (.B1(_1641_),
    .Y(_1642_),
    .A1(_1637_),
    .A2(_1640_));
 sg13g2_inv_1 _3196_ (.Y(_0184_),
    .A(net545));
 sg13g2_nand2b_1 _3197_ (.Y(_1643_),
    .B(\s0.data_out[6][7] ),
    .A_N(net1021));
 sg13g2_a21oi_1 _3198_ (.A1(_1552_),
    .A2(_1643_),
    .Y(_1644_),
    .B1(net1018));
 sg13g2_nor2b_1 _3199_ (.A(net1006),
    .B_N(net1047),
    .Y(_1645_));
 sg13g2_a21oi_1 _3200_ (.A1(net1006),
    .A2(\s0.data_out[6][7] ),
    .Y(_1646_),
    .B1(_1645_));
 sg13g2_o21ai_1 _3201_ (.B1(net1329),
    .Y(_1647_),
    .A1(net917),
    .A2(_1646_));
 sg13g2_or2_1 _3202_ (.X(_1648_),
    .B(net517),
    .A(net1329));
 sg13g2_o21ai_1 _3203_ (.B1(_1648_),
    .Y(_1649_),
    .A1(_1644_),
    .A2(_1647_));
 sg13g2_inv_1 _3204_ (.Y(_0185_),
    .A(net518));
 sg13g2_nand2_1 _3205_ (.Y(_1650_),
    .A(net1011),
    .B(net484));
 sg13g2_o21ai_1 _3206_ (.B1(_1650_),
    .Y(_1651_),
    .A1(net1008),
    .A2(_2491_));
 sg13g2_a21oi_1 _3207_ (.A1(net1001),
    .A2(_1651_),
    .Y(_1652_),
    .B1(_1611_));
 sg13g2_o21ai_1 _3208_ (.B1(_1609_),
    .Y(_1653_),
    .A1(net917),
    .A2(_1652_));
 sg13g2_nand2_1 _3209_ (.Y(_1654_),
    .A(net1008),
    .B(net537));
 sg13g2_mux2_1 _3210_ (.A0(\s0.data_out[7][1] ),
    .A1(\s0.data_out[6][1] ),
    .S(net1008),
    .X(_1655_));
 sg13g2_a21oi_1 _3211_ (.A1(net1001),
    .A2(_1655_),
    .Y(_1656_),
    .B1(_1604_));
 sg13g2_nand2b_1 _3212_ (.Y(_1657_),
    .B(net1012),
    .A_N(_1656_));
 sg13g2_nand3_1 _3213_ (.B(_1602_),
    .C(_1657_),
    .A(net1278),
    .Y(_1658_));
 sg13g2_mux2_1 _3214_ (.A0(\s0.data_out[7][0] ),
    .A1(\s0.data_out[6][0] ),
    .S(net1011),
    .X(_1659_));
 sg13g2_a21oi_1 _3215_ (.A1(net1001),
    .A2(_1659_),
    .Y(_1660_),
    .B1(_1597_));
 sg13g2_o21ai_1 _3216_ (.B1(_1595_),
    .Y(_1661_),
    .A1(net917),
    .A2(_1660_));
 sg13g2_nor2b_1 _3217_ (.A(net1282),
    .B_N(_1661_),
    .Y(_1662_));
 sg13g2_a21oi_1 _3218_ (.A1(_1602_),
    .A2(_1657_),
    .Y(_1663_),
    .B1(net1278));
 sg13g2_a221oi_1 _3219_ (.B2(_1662_),
    .C1(_1663_),
    .B1(_1658_),
    .A1(net1212),
    .Y(_1664_),
    .A2(_1653_));
 sg13g2_mux2_1 _3220_ (.A0(\s0.data_out[7][3] ),
    .A1(\s0.data_out[6][3] ),
    .S(net1011),
    .X(_1665_));
 sg13g2_a21o_1 _3221_ (.A2(_1665_),
    .A1(net1002),
    .B1(_1617_),
    .X(_1666_));
 sg13g2_a21oi_1 _3222_ (.A1(net1014),
    .A2(_1666_),
    .Y(_1667_),
    .B1(_1616_));
 sg13g2_nand2_1 _3223_ (.Y(_1668_),
    .A(net1264),
    .B(_1667_));
 sg13g2_o21ai_1 _3224_ (.B1(_1668_),
    .Y(_1669_),
    .A1(net1212),
    .A2(_1653_));
 sg13g2_mux2_1 _3225_ (.A0(\s0.data_out[7][4] ),
    .A1(\s0.data_out[6][4] ),
    .S(net1009),
    .X(_1670_));
 sg13g2_a21o_1 _3226_ (.A2(_1670_),
    .A1(net1005),
    .B1(_1624_),
    .X(_1671_));
 sg13g2_a21oi_1 _3227_ (.A1(net1015),
    .A2(_1671_),
    .Y(_1672_),
    .B1(_1623_));
 sg13g2_nand2_1 _3228_ (.Y(_1673_),
    .A(net1009),
    .B(net539));
 sg13g2_mux2_1 _3229_ (.A0(\s0.data_out[7][5] ),
    .A1(\s0.data_out[6][5] ),
    .S(net1010),
    .X(_1674_));
 sg13g2_a21o_1 _3230_ (.A2(_1674_),
    .A1(net1005),
    .B1(_1631_),
    .X(_1675_));
 sg13g2_a21oi_1 _3231_ (.A1(net1015),
    .A2(_1675_),
    .Y(_1676_),
    .B1(_1630_));
 sg13g2_a22oi_1 _3232_ (.Y(_1677_),
    .B1(_1676_),
    .B2(net1250),
    .A2(_1672_),
    .A1(net1258));
 sg13g2_nor2_1 _3233_ (.A(net1250),
    .B(_1676_),
    .Y(_1678_));
 sg13g2_nor2_1 _3234_ (.A(net1258),
    .B(_1672_),
    .Y(_1679_));
 sg13g2_nor2_1 _3235_ (.A(net1264),
    .B(_1667_),
    .Y(_1680_));
 sg13g2_nor3_1 _3236_ (.A(_1678_),
    .B(_1679_),
    .C(_1680_),
    .Y(_1681_));
 sg13g2_nand2_1 _3237_ (.Y(_1682_),
    .A(_1677_),
    .B(_1681_));
 sg13g2_nand2_1 _3238_ (.Y(_1683_),
    .A(net1009),
    .B(net519));
 sg13g2_mux2_1 _3239_ (.A0(\s0.data_out[7][7] ),
    .A1(\s0.data_out[6][7] ),
    .S(net1010),
    .X(_1684_));
 sg13g2_a21o_1 _3240_ (.A2(_1684_),
    .A1(net1006),
    .B1(_1645_),
    .X(_1685_));
 sg13g2_a21oi_1 _3241_ (.A1(net1018),
    .A2(_1685_),
    .Y(_1686_),
    .B1(_1644_));
 sg13g2_nand2_1 _3242_ (.Y(_1687_),
    .A(net1009),
    .B(net557));
 sg13g2_mux2_1 _3243_ (.A0(\s0.data_out[7][6] ),
    .A1(\s0.data_out[6][6] ),
    .S(net1010),
    .X(_1688_));
 sg13g2_a21o_1 _3244_ (.A2(_1688_),
    .A1(net1006),
    .B1(_1638_),
    .X(_1689_));
 sg13g2_a21oi_1 _3245_ (.A1(net1015),
    .A2(_1689_),
    .Y(_1690_),
    .B1(_1637_));
 sg13g2_a22oi_1 _3246_ (.Y(_1691_),
    .B1(_1690_),
    .B2(net1244),
    .A2(_1686_),
    .A1(net1235));
 sg13g2_or2_1 _3247_ (.X(_1692_),
    .B(_1690_),
    .A(net1244));
 sg13g2_nor2_1 _3248_ (.A(net1235),
    .B(_1686_),
    .Y(_1693_));
 sg13g2_or2_1 _3249_ (.X(_1694_),
    .B(_1686_),
    .A(net1238));
 sg13g2_and3_1 _3250_ (.X(_1695_),
    .A(_1691_),
    .B(_1692_),
    .C(_1694_));
 sg13g2_o21ai_1 _3251_ (.B1(_1695_),
    .Y(_1696_),
    .A1(_1664_),
    .A2(_1669_));
 sg13g2_nor2_1 _3252_ (.A(_1677_),
    .B(_1678_),
    .Y(_1697_));
 sg13g2_o21ai_1 _3253_ (.B1(_1592_),
    .Y(_1698_),
    .A1(_1691_),
    .A2(_1693_));
 sg13g2_a21oi_1 _3254_ (.A1(_1695_),
    .A2(_1697_),
    .Y(_1699_),
    .B1(_1698_));
 sg13g2_o21ai_1 _3255_ (.B1(_1699_),
    .Y(_1700_),
    .A1(_1682_),
    .A2(_1696_));
 sg13g2_nor2_1 _3256_ (.A(net313),
    .B(net1209),
    .Y(_1701_));
 sg13g2_and2_1 _3257_ (.A(_1700_),
    .B(_1701_),
    .X(_0186_));
 sg13g2_and2_1 _3258_ (.A(net1325),
    .B(net309),
    .X(_0187_));
 sg13g2_o21ai_1 _3259_ (.B1(net1004),
    .Y(_1702_),
    .A1(net1230),
    .A2(net995));
 sg13g2_nor2b_1 _3260_ (.A(net1230),
    .B_N(net999),
    .Y(_1703_));
 sg13g2_nor2_1 _3261_ (.A(_1702_),
    .B(_1703_),
    .Y(_1704_));
 sg13g2_inv_1 _3262_ (.Y(_1705_),
    .A(_1704_));
 sg13g2_o21ai_1 _3263_ (.B1(_1705_),
    .Y(_1706_),
    .A1(net1004),
    .A2(_1585_));
 sg13g2_or2_1 _3264_ (.X(_1707_),
    .B(net999),
    .A(net383));
 sg13g2_o21ai_1 _3265_ (.B1(_2469_),
    .Y(_1708_),
    .A1(net383),
    .A2(net1009));
 sg13g2_o21ai_1 _3266_ (.B1(_1708_),
    .Y(_1709_),
    .A1(net995),
    .A2(_1702_));
 sg13g2_a21oi_1 _3267_ (.A1(_1704_),
    .A2(_1707_),
    .Y(_1710_),
    .B1(_1709_));
 sg13g2_o21ai_1 _3268_ (.B1(net1325),
    .Y(_1711_),
    .A1(net465),
    .A2(_1706_));
 sg13g2_nor2_1 _3269_ (.A(_1710_),
    .B(_1711_),
    .Y(_0188_));
 sg13g2_nor2_1 _3270_ (.A(net1220),
    .B(_1706_),
    .Y(_0189_));
 sg13g2_mux2_1 _3271_ (.A0(\s0.data_out[5][0] ),
    .A1(\s0.data_out[6][0] ),
    .S(net1008),
    .X(_1712_));
 sg13g2_nand2_1 _3272_ (.Y(_1713_),
    .A(net916),
    .B(_1712_));
 sg13g2_and2_1 _3273_ (.A(net991),
    .B(\s0.data_out[5][0] ),
    .X(_1714_));
 sg13g2_nor2b_1 _3274_ (.A(net991),
    .B_N(net1074),
    .Y(_1715_));
 sg13g2_o21ai_1 _3275_ (.B1(net1000),
    .Y(_1716_),
    .A1(_1714_),
    .A2(_1715_));
 sg13g2_nand3_1 _3276_ (.B(_1713_),
    .C(_1716_),
    .A(net1324),
    .Y(_1717_));
 sg13g2_o21ai_1 _3277_ (.B1(_1717_),
    .Y(_1718_),
    .A1(net1326),
    .A2(net412));
 sg13g2_inv_1 _3278_ (.Y(_0190_),
    .A(_1718_));
 sg13g2_nand2b_1 _3279_ (.Y(_1719_),
    .B(net463),
    .A_N(net1008));
 sg13g2_a21oi_1 _3280_ (.A1(_1654_),
    .A2(_1719_),
    .Y(_1720_),
    .B1(net1000));
 sg13g2_nor2b_1 _3281_ (.A(net992),
    .B_N(net1070),
    .Y(_1721_));
 sg13g2_a21oi_1 _3282_ (.A1(net991),
    .A2(net463),
    .Y(_1722_),
    .B1(_1721_));
 sg13g2_o21ai_1 _3283_ (.B1(net1324),
    .Y(_1723_),
    .A1(net916),
    .A2(_1722_));
 sg13g2_or2_1 _3284_ (.X(_1724_),
    .B(net537),
    .A(net1324));
 sg13g2_o21ai_1 _3285_ (.B1(_1724_),
    .Y(_1725_),
    .A1(_1720_),
    .A2(_1723_));
 sg13g2_inv_1 _3286_ (.Y(_0191_),
    .A(_1725_));
 sg13g2_nand2b_1 _3287_ (.Y(_1726_),
    .B(\s0.data_out[5][2] ),
    .A_N(net1008));
 sg13g2_a21oi_1 _3288_ (.A1(_1650_),
    .A2(_1726_),
    .Y(_1727_),
    .B1(net1000));
 sg13g2_nor2b_1 _3289_ (.A(net991),
    .B_N(net1066),
    .Y(_1728_));
 sg13g2_a21oi_1 _3290_ (.A1(net991),
    .A2(\s0.data_out[5][2] ),
    .Y(_1729_),
    .B1(_1728_));
 sg13g2_o21ai_1 _3291_ (.B1(net1326),
    .Y(_1730_),
    .A1(net916),
    .A2(_1729_));
 sg13g2_or2_1 _3292_ (.X(_1731_),
    .B(net484),
    .A(net1324));
 sg13g2_o21ai_1 _3293_ (.B1(_1731_),
    .Y(_1732_),
    .A1(_1727_),
    .A2(_1730_));
 sg13g2_inv_1 _3294_ (.Y(_0192_),
    .A(net485));
 sg13g2_mux2_1 _3295_ (.A0(\s0.data_out[5][3] ),
    .A1(\s0.data_out[6][3] ),
    .S(net1008),
    .X(_1733_));
 sg13g2_nand2_1 _3296_ (.Y(_1734_),
    .A(net916),
    .B(_1733_));
 sg13g2_and2_1 _3297_ (.A(net992),
    .B(\s0.data_out[5][3] ),
    .X(_1735_));
 sg13g2_nor2b_1 _3298_ (.A(net992),
    .B_N(net1062),
    .Y(_1736_));
 sg13g2_o21ai_1 _3299_ (.B1(net1000),
    .Y(_1737_),
    .A1(_1735_),
    .A2(_1736_));
 sg13g2_nand3_1 _3300_ (.B(_1734_),
    .C(_1737_),
    .A(net1324),
    .Y(_1738_));
 sg13g2_o21ai_1 _3301_ (.B1(_1738_),
    .Y(_1739_),
    .A1(net1324),
    .A2(net454));
 sg13g2_inv_1 _3302_ (.Y(_0193_),
    .A(_1739_));
 sg13g2_mux2_1 _3303_ (.A0(\s0.data_out[5][4] ),
    .A1(\s0.data_out[6][4] ),
    .S(net1008),
    .X(_1740_));
 sg13g2_nand2_1 _3304_ (.Y(_1741_),
    .A(net916),
    .B(_1740_));
 sg13g2_and2_1 _3305_ (.A(net992),
    .B(\s0.data_out[5][4] ),
    .X(_1742_));
 sg13g2_nor2b_1 _3306_ (.A(net992),
    .B_N(net1059),
    .Y(_1743_));
 sg13g2_o21ai_1 _3307_ (.B1(net1000),
    .Y(_1744_),
    .A1(_1742_),
    .A2(_1743_));
 sg13g2_nand3_1 _3308_ (.B(_1741_),
    .C(_1744_),
    .A(net1326),
    .Y(_1745_));
 sg13g2_o21ai_1 _3309_ (.B1(_1745_),
    .Y(_1746_),
    .A1(net1324),
    .A2(net423));
 sg13g2_inv_1 _3310_ (.Y(_0194_),
    .A(_1746_));
 sg13g2_nand2b_1 _3311_ (.Y(_1747_),
    .B(net352),
    .A_N(net1009));
 sg13g2_a21oi_1 _3312_ (.A1(_1673_),
    .A2(_1747_),
    .Y(_1748_),
    .B1(net1004));
 sg13g2_nor2b_1 _3313_ (.A(net995),
    .B_N(net1055),
    .Y(_1749_));
 sg13g2_a21oi_1 _3314_ (.A1(net995),
    .A2(net352),
    .Y(_1750_),
    .B1(_1749_));
 sg13g2_o21ai_1 _3315_ (.B1(net1325),
    .Y(_1751_),
    .A1(net916),
    .A2(_1750_));
 sg13g2_or2_1 _3316_ (.X(_1752_),
    .B(net539),
    .A(net1325));
 sg13g2_o21ai_1 _3317_ (.B1(_1752_),
    .Y(_1753_),
    .A1(_1748_),
    .A2(_1751_));
 sg13g2_inv_1 _3318_ (.Y(_0195_),
    .A(_1753_));
 sg13g2_nand2b_1 _3319_ (.Y(_1754_),
    .B(net538),
    .A_N(net1009));
 sg13g2_a21oi_1 _3320_ (.A1(_1687_),
    .A2(_1754_),
    .Y(_1755_),
    .B1(net1004));
 sg13g2_nor2b_1 _3321_ (.A(net996),
    .B_N(net1051),
    .Y(_1756_));
 sg13g2_a21oi_1 _3322_ (.A1(net996),
    .A2(net538),
    .Y(_1757_),
    .B1(_1756_));
 sg13g2_o21ai_1 _3323_ (.B1(net1325),
    .Y(_1758_),
    .A1(net916),
    .A2(_1757_));
 sg13g2_or2_1 _3324_ (.X(_1759_),
    .B(net557),
    .A(net1325));
 sg13g2_o21ai_1 _3325_ (.B1(_1759_),
    .Y(_1760_),
    .A1(_1755_),
    .A2(_1758_));
 sg13g2_inv_1 _3326_ (.Y(_0196_),
    .A(_1760_));
 sg13g2_nand2b_1 _3327_ (.Y(_1761_),
    .B(\s0.data_out[5][7] ),
    .A_N(net1009));
 sg13g2_a21oi_1 _3328_ (.A1(_1683_),
    .A2(_1761_),
    .Y(_1762_),
    .B1(net1004));
 sg13g2_nor2b_1 _3329_ (.A(net996),
    .B_N(net1047),
    .Y(_1763_));
 sg13g2_a21oi_1 _3330_ (.A1(net995),
    .A2(\s0.data_out[5][7] ),
    .Y(_1764_),
    .B1(_1763_));
 sg13g2_o21ai_1 _3331_ (.B1(net1325),
    .Y(_1765_),
    .A1(net916),
    .A2(_1764_));
 sg13g2_or2_1 _3332_ (.X(_1766_),
    .B(net519),
    .A(net1325));
 sg13g2_o21ai_1 _3333_ (.B1(_1766_),
    .Y(_1767_),
    .A1(_1762_),
    .A2(_1765_));
 sg13g2_inv_1 _3334_ (.Y(_0197_),
    .A(net520));
 sg13g2_nand2_1 _3335_ (.Y(_1768_),
    .A(net997),
    .B(net581));
 sg13g2_mux2_1 _3336_ (.A0(\s0.data_out[6][2] ),
    .A1(\s0.data_out[5][2] ),
    .S(net999),
    .X(_1769_));
 sg13g2_a21o_1 _3337_ (.A2(_1769_),
    .A1(net991),
    .B1(_1728_),
    .X(_1770_));
 sg13g2_a21oi_1 _3338_ (.A1(net1000),
    .A2(_1770_),
    .Y(_1771_),
    .B1(_1727_));
 sg13g2_or2_1 _3339_ (.X(_1772_),
    .B(_1771_),
    .A(net1271));
 sg13g2_mux2_1 _3340_ (.A0(\s0.data_out[6][1] ),
    .A1(\s0.data_out[5][1] ),
    .S(net997),
    .X(_1773_));
 sg13g2_a21o_1 _3341_ (.A2(_1773_),
    .A1(net991),
    .B1(_1721_),
    .X(_1774_));
 sg13g2_a21oi_1 _3342_ (.A1(net1000),
    .A2(_1774_),
    .Y(_1775_),
    .B1(_1720_));
 sg13g2_mux2_1 _3343_ (.A0(\s0.data_out[6][0] ),
    .A1(\s0.data_out[5][0] ),
    .S(net997),
    .X(_1776_));
 sg13g2_a21oi_1 _3344_ (.A1(net991),
    .A2(_1776_),
    .Y(_1777_),
    .B1(_1715_));
 sg13g2_nand2b_1 _3345_ (.Y(_1778_),
    .B(net1000),
    .A_N(_1777_));
 sg13g2_o21ai_1 _3346_ (.B1(_1772_),
    .Y(_1779_),
    .A1(net1277),
    .A2(_1775_));
 sg13g2_a221oi_1 _3347_ (.B2(_1713_),
    .C1(net1282),
    .B1(_1778_),
    .A1(net1277),
    .Y(_1780_),
    .A2(_1775_));
 sg13g2_mux2_1 _3348_ (.A0(\s0.data_out[6][3] ),
    .A1(\s0.data_out[5][3] ),
    .S(net999),
    .X(_1781_));
 sg13g2_a21oi_1 _3349_ (.A1(net992),
    .A2(_1781_),
    .Y(_1782_),
    .B1(_1736_));
 sg13g2_nand2b_1 _3350_ (.Y(_1783_),
    .B(net1003),
    .A_N(_1782_));
 sg13g2_and2_1 _3351_ (.A(_1734_),
    .B(_1783_),
    .X(_1784_));
 sg13g2_a22oi_1 _3352_ (.Y(_1785_),
    .B1(_1784_),
    .B2(net1264),
    .A2(_1771_),
    .A1(net1271));
 sg13g2_o21ai_1 _3353_ (.B1(_1785_),
    .Y(_1786_),
    .A1(_1779_),
    .A2(_1780_));
 sg13g2_nand2_1 _3354_ (.Y(_1787_),
    .A(net998),
    .B(net569));
 sg13g2_mux2_1 _3355_ (.A0(\s0.data_out[6][7] ),
    .A1(\s0.data_out[5][7] ),
    .S(net998),
    .X(_1788_));
 sg13g2_a21o_1 _3356_ (.A2(_1788_),
    .A1(net995),
    .B1(_1763_),
    .X(_1789_));
 sg13g2_a21oi_1 _3357_ (.A1(net1007),
    .A2(_1789_),
    .Y(_1790_),
    .B1(_1762_));
 sg13g2_nand2_1 _3358_ (.Y(_1791_),
    .A(net998),
    .B(net538));
 sg13g2_mux2_1 _3359_ (.A0(\s0.data_out[6][6] ),
    .A1(\s0.data_out[5][6] ),
    .S(net999),
    .X(_1792_));
 sg13g2_a21o_1 _3360_ (.A2(_1792_),
    .A1(net995),
    .B1(_1756_),
    .X(_1793_));
 sg13g2_a21oi_1 _3361_ (.A1(net1004),
    .A2(_1793_),
    .Y(_1794_),
    .B1(_1755_));
 sg13g2_a22oi_1 _3362_ (.Y(_1795_),
    .B1(_1794_),
    .B2(net1244),
    .A2(_1790_),
    .A1(net1235));
 sg13g2_nor2_1 _3363_ (.A(net1244),
    .B(_1794_),
    .Y(_1796_));
 sg13g2_or2_1 _3364_ (.X(_1797_),
    .B(_1790_),
    .A(net1235));
 sg13g2_nand3b_1 _3365_ (.B(_1797_),
    .C(_1795_),
    .Y(_1798_),
    .A_N(_1796_));
 sg13g2_mux2_1 _3366_ (.A0(\s0.data_out[6][5] ),
    .A1(\s0.data_out[5][5] ),
    .S(net998),
    .X(_1799_));
 sg13g2_a21o_1 _3367_ (.A2(_1799_),
    .A1(net995),
    .B1(_1749_),
    .X(_1800_));
 sg13g2_a21oi_1 _3368_ (.A1(net1004),
    .A2(_1800_),
    .Y(_1801_),
    .B1(_1748_));
 sg13g2_nand2_1 _3369_ (.Y(_1802_),
    .A(net1250),
    .B(_1801_));
 sg13g2_o21ai_1 _3370_ (.B1(_1802_),
    .Y(_1803_),
    .A1(net1264),
    .A2(_1784_));
 sg13g2_mux2_1 _3371_ (.A0(\s0.data_out[6][4] ),
    .A1(\s0.data_out[5][4] ),
    .S(net999),
    .X(_1804_));
 sg13g2_a21oi_1 _3372_ (.A1(net992),
    .A2(_1804_),
    .Y(_1805_),
    .B1(_1743_));
 sg13g2_nand2b_1 _3373_ (.Y(_1806_),
    .B(net1003),
    .A_N(_1805_));
 sg13g2_a21o_1 _3374_ (.A2(_1806_),
    .A1(_1741_),
    .B1(net1258),
    .X(_1807_));
 sg13g2_nand3_1 _3375_ (.B(_1741_),
    .C(_1806_),
    .A(net1258),
    .Y(_1808_));
 sg13g2_nor2_1 _3376_ (.A(net1250),
    .B(_1801_),
    .Y(_1809_));
 sg13g2_nor3_1 _3377_ (.A(_1798_),
    .B(_1803_),
    .C(_1809_),
    .Y(_1810_));
 sg13g2_nand4_1 _3378_ (.B(_1807_),
    .C(_1808_),
    .A(_1786_),
    .Y(_1811_),
    .D(_1810_));
 sg13g2_o21ai_1 _3379_ (.B1(_1802_),
    .Y(_1812_),
    .A1(_1808_),
    .A2(_1809_));
 sg13g2_nor2b_1 _3380_ (.A(_1798_),
    .B_N(_1812_),
    .Y(_1813_));
 sg13g2_nor2b_1 _3381_ (.A(_1795_),
    .B_N(_1797_),
    .Y(_1814_));
 sg13g2_nor3_1 _3382_ (.A(_1706_),
    .B(_1813_),
    .C(_1814_),
    .Y(_1815_));
 sg13g2_or2_1 _3383_ (.X(_1816_),
    .B(net1209),
    .A(net309));
 sg13g2_a21oi_1 _3384_ (.A1(_1811_),
    .A2(_1815_),
    .Y(_0198_),
    .B1(_1816_));
 sg13g2_and2_1 _3385_ (.A(net1313),
    .B(net318),
    .X(_0199_));
 sg13g2_o21ai_1 _3386_ (.B1(net994),
    .Y(_1817_),
    .A1(net1226),
    .A2(net984));
 sg13g2_nor2b_1 _3387_ (.A(net1226),
    .B_N(net989),
    .Y(_1818_));
 sg13g2_nor2_1 _3388_ (.A(_1817_),
    .B(_1818_),
    .Y(_1819_));
 sg13g2_nor2_1 _3389_ (.A(net994),
    .B(_1703_),
    .Y(_1820_));
 sg13g2_or2_1 _3390_ (.X(_1821_),
    .B(_1820_),
    .A(_1819_));
 sg13g2_or2_1 _3391_ (.X(_1822_),
    .B(net989),
    .A(net353));
 sg13g2_o21ai_1 _3392_ (.B1(net915),
    .Y(_1823_),
    .A1(net353),
    .A2(net998));
 sg13g2_o21ai_1 _3393_ (.B1(_1823_),
    .Y(_1824_),
    .A1(net985),
    .A2(_1817_));
 sg13g2_a21oi_1 _3394_ (.A1(_1819_),
    .A2(_1822_),
    .Y(_1825_),
    .B1(_1824_));
 sg13g2_o21ai_1 _3395_ (.B1(net1313),
    .Y(_1826_),
    .A1(net383),
    .A2(_1821_));
 sg13g2_nor2_1 _3396_ (.A(_1825_),
    .B(_1826_),
    .Y(_0200_));
 sg13g2_nor2_1 _3397_ (.A(net1219),
    .B(_1821_),
    .Y(_0201_));
 sg13g2_mux2_1 _3398_ (.A0(\s0.data_out[4][0] ),
    .A1(\s0.data_out[5][0] ),
    .S(net997),
    .X(_1827_));
 sg13g2_nand2_1 _3399_ (.Y(_1828_),
    .A(net915),
    .B(_1827_));
 sg13g2_and2_1 _3400_ (.A(net981),
    .B(\s0.data_out[4][0] ),
    .X(_1829_));
 sg13g2_nor2b_1 _3401_ (.A(net981),
    .B_N(net1074),
    .Y(_1830_));
 sg13g2_o21ai_1 _3402_ (.B1(net990),
    .Y(_1831_),
    .A1(_1829_),
    .A2(_1830_));
 sg13g2_nand3_1 _3403_ (.B(_1828_),
    .C(_1831_),
    .A(net1311),
    .Y(_1832_));
 sg13g2_o21ai_1 _3404_ (.B1(_1832_),
    .Y(_1833_),
    .A1(net1311),
    .A2(net432));
 sg13g2_inv_1 _3405_ (.Y(_0202_),
    .A(_1833_));
 sg13g2_mux2_1 _3406_ (.A0(\s0.data_out[4][1] ),
    .A1(\s0.data_out[5][1] ),
    .S(net997),
    .X(_1834_));
 sg13g2_nand2_1 _3407_ (.Y(_1835_),
    .A(net915),
    .B(_1834_));
 sg13g2_and2_1 _3408_ (.A(net982),
    .B(\s0.data_out[4][1] ),
    .X(_1836_));
 sg13g2_nor2b_1 _3409_ (.A(net981),
    .B_N(net1070),
    .Y(_1837_));
 sg13g2_o21ai_1 _3410_ (.B1(net990),
    .Y(_1838_),
    .A1(_1836_),
    .A2(_1837_));
 sg13g2_nand3_1 _3411_ (.B(_1835_),
    .C(_1838_),
    .A(net1311),
    .Y(_1839_));
 sg13g2_o21ai_1 _3412_ (.B1(_1839_),
    .Y(_1840_),
    .A1(net1311),
    .A2(net463));
 sg13g2_inv_1 _3413_ (.Y(_0203_),
    .A(_1840_));
 sg13g2_nand2b_1 _3414_ (.Y(_1841_),
    .B(net533),
    .A_N(net997));
 sg13g2_a21oi_1 _3415_ (.A1(_1768_),
    .A2(_1841_),
    .Y(_1842_),
    .B1(net990));
 sg13g2_nor2b_1 _3416_ (.A(net981),
    .B_N(net1066),
    .Y(_1843_));
 sg13g2_a21oi_1 _3417_ (.A1(net981),
    .A2(net533),
    .Y(_1844_),
    .B1(_1843_));
 sg13g2_o21ai_1 _3418_ (.B1(net1311),
    .Y(_1845_),
    .A1(net915),
    .A2(_1844_));
 sg13g2_or2_1 _3419_ (.X(_1846_),
    .B(net581),
    .A(net1311));
 sg13g2_o21ai_1 _3420_ (.B1(_1846_),
    .Y(_1847_),
    .A1(_1842_),
    .A2(_1845_));
 sg13g2_inv_1 _3421_ (.Y(_0204_),
    .A(_1847_));
 sg13g2_mux2_1 _3422_ (.A0(\s0.data_out[4][3] ),
    .A1(\s0.data_out[5][3] ),
    .S(net997),
    .X(_1848_));
 sg13g2_nand2_1 _3423_ (.Y(_1849_),
    .A(net915),
    .B(_1848_));
 sg13g2_and2_1 _3424_ (.A(net982),
    .B(\s0.data_out[4][3] ),
    .X(_1850_));
 sg13g2_nor2b_1 _3425_ (.A(net982),
    .B_N(net1062),
    .Y(_1851_));
 sg13g2_o21ai_1 _3426_ (.B1(net990),
    .Y(_1852_),
    .A1(_1850_),
    .A2(_1851_));
 sg13g2_nand3_1 _3427_ (.B(_1849_),
    .C(_1852_),
    .A(net1311),
    .Y(_1853_));
 sg13g2_o21ai_1 _3428_ (.B1(_1853_),
    .Y(_1854_),
    .A1(net1311),
    .A2(net415));
 sg13g2_inv_1 _3429_ (.Y(_0205_),
    .A(_1854_));
 sg13g2_mux2_1 _3430_ (.A0(\s0.data_out[4][4] ),
    .A1(\s0.data_out[5][4] ),
    .S(net997),
    .X(_1855_));
 sg13g2_nand2_1 _3431_ (.Y(_1856_),
    .A(net915),
    .B(_1855_));
 sg13g2_and2_1 _3432_ (.A(net982),
    .B(\s0.data_out[4][4] ),
    .X(_1857_));
 sg13g2_nor2b_1 _3433_ (.A(net982),
    .B_N(net1058),
    .Y(_1858_));
 sg13g2_o21ai_1 _3434_ (.B1(net993),
    .Y(_1859_),
    .A1(_1857_),
    .A2(_1858_));
 sg13g2_nand3_1 _3435_ (.B(_1856_),
    .C(_1859_),
    .A(net1312),
    .Y(_1860_));
 sg13g2_o21ai_1 _3436_ (.B1(_1860_),
    .Y(_1861_),
    .A1(net1315),
    .A2(net402));
 sg13g2_inv_1 _3437_ (.Y(_0206_),
    .A(_1861_));
 sg13g2_mux2_1 _3438_ (.A0(\s0.data_out[4][5] ),
    .A1(\s0.data_out[5][5] ),
    .S(net998),
    .X(_1862_));
 sg13g2_nand2_1 _3439_ (.Y(_1863_),
    .A(net915),
    .B(_1862_));
 sg13g2_and2_1 _3440_ (.A(net984),
    .B(\s0.data_out[4][5] ),
    .X(_1864_));
 sg13g2_nor2b_1 _3441_ (.A(net984),
    .B_N(net1054),
    .Y(_1865_));
 sg13g2_o21ai_1 _3442_ (.B1(net994),
    .Y(_1866_),
    .A1(_1864_),
    .A2(_1865_));
 sg13g2_nand3_1 _3443_ (.B(_1863_),
    .C(_1866_),
    .A(net1314),
    .Y(_1867_));
 sg13g2_o21ai_1 _3444_ (.B1(_1867_),
    .Y(_1868_),
    .A1(net1314),
    .A2(net352));
 sg13g2_inv_1 _3445_ (.Y(_0207_),
    .A(_1868_));
 sg13g2_nand2b_1 _3446_ (.Y(_1869_),
    .B(net511),
    .A_N(net998));
 sg13g2_a21oi_1 _3447_ (.A1(_1791_),
    .A2(_1869_),
    .Y(_1870_),
    .B1(net994));
 sg13g2_nor2b_1 _3448_ (.A(net985),
    .B_N(net1050),
    .Y(_1871_));
 sg13g2_a21oi_1 _3449_ (.A1(net985),
    .A2(net511),
    .Y(_1872_),
    .B1(_1871_));
 sg13g2_o21ai_1 _3450_ (.B1(net1314),
    .Y(_1873_),
    .A1(_2470_),
    .A2(_1872_));
 sg13g2_or2_1 _3451_ (.X(_1874_),
    .B(net538),
    .A(net1313));
 sg13g2_o21ai_1 _3452_ (.B1(_1874_),
    .Y(_1875_),
    .A1(_1870_),
    .A2(_1873_));
 sg13g2_inv_1 _3453_ (.Y(_0208_),
    .A(_1875_));
 sg13g2_nand2b_1 _3454_ (.Y(_1876_),
    .B(net535),
    .A_N(net998));
 sg13g2_a21oi_1 _3455_ (.A1(_1787_),
    .A2(_1876_),
    .Y(_1877_),
    .B1(net994));
 sg13g2_nor2b_1 _3456_ (.A(net984),
    .B_N(net1046),
    .Y(_1878_));
 sg13g2_a21oi_1 _3457_ (.A1(net984),
    .A2(net535),
    .Y(_1879_),
    .B1(_1878_));
 sg13g2_o21ai_1 _3458_ (.B1(net1314),
    .Y(_1880_),
    .A1(net915),
    .A2(_1879_));
 sg13g2_or2_1 _3459_ (.X(_1881_),
    .B(net569),
    .A(net1314));
 sg13g2_o21ai_1 _3460_ (.B1(_1881_),
    .Y(_1882_),
    .A1(_1877_),
    .A2(_1880_));
 sg13g2_inv_1 _3461_ (.Y(_0209_),
    .A(_1882_));
 sg13g2_nand2_1 _3462_ (.Y(_1883_),
    .A(net987),
    .B(net533));
 sg13g2_mux2_1 _3463_ (.A0(\s0.data_out[5][2] ),
    .A1(\s0.data_out[4][2] ),
    .S(net987),
    .X(_1884_));
 sg13g2_a21o_1 _3464_ (.A2(_1884_),
    .A1(net981),
    .B1(_1843_),
    .X(_1885_));
 sg13g2_a21oi_1 _3465_ (.A1(net990),
    .A2(_1885_),
    .Y(_1886_),
    .B1(_1842_));
 sg13g2_or2_1 _3466_ (.X(_1887_),
    .B(_1886_),
    .A(net1271));
 sg13g2_mux2_1 _3467_ (.A0(\s0.data_out[5][1] ),
    .A1(\s0.data_out[4][1] ),
    .S(net987),
    .X(_1888_));
 sg13g2_a21oi_1 _3468_ (.A1(net981),
    .A2(_1888_),
    .Y(_1889_),
    .B1(_1837_));
 sg13g2_nand2b_1 _3469_ (.Y(_1890_),
    .B(net990),
    .A_N(_1889_));
 sg13g2_and2_1 _3470_ (.A(_1835_),
    .B(_1890_),
    .X(_1891_));
 sg13g2_mux2_1 _3471_ (.A0(\s0.data_out[5][0] ),
    .A1(\s0.data_out[4][0] ),
    .S(net989),
    .X(_1892_));
 sg13g2_a21oi_1 _3472_ (.A1(net981),
    .A2(_1892_),
    .Y(_1893_),
    .B1(_1830_));
 sg13g2_nand2b_1 _3473_ (.Y(_1894_),
    .B(net990),
    .A_N(_1893_));
 sg13g2_a221oi_1 _3474_ (.B2(_1828_),
    .C1(net1282),
    .B1(_1894_),
    .A1(net1277),
    .Y(_1895_),
    .A2(_1891_));
 sg13g2_o21ai_1 _3475_ (.B1(_1887_),
    .Y(_1896_),
    .A1(net1280),
    .A2(_1891_));
 sg13g2_mux2_1 _3476_ (.A0(\s0.data_out[5][3] ),
    .A1(\s0.data_out[4][3] ),
    .S(net989),
    .X(_1897_));
 sg13g2_a21oi_1 _3477_ (.A1(net982),
    .A2(_1897_),
    .Y(_1898_),
    .B1(_1851_));
 sg13g2_nand2b_1 _3478_ (.Y(_1899_),
    .B(net990),
    .A_N(_1898_));
 sg13g2_and2_1 _3479_ (.A(_1849_),
    .B(_1899_),
    .X(_1900_));
 sg13g2_a22oi_1 _3480_ (.Y(_1901_),
    .B1(_1900_),
    .B2(net1267),
    .A2(_1886_),
    .A1(net1271));
 sg13g2_o21ai_1 _3481_ (.B1(_1901_),
    .Y(_1902_),
    .A1(_1895_),
    .A2(_1896_));
 sg13g2_nand2_1 _3482_ (.Y(_1903_),
    .A(net988),
    .B(net535));
 sg13g2_mux2_1 _3483_ (.A0(\s0.data_out[5][7] ),
    .A1(\s0.data_out[4][7] ),
    .S(net988),
    .X(_1904_));
 sg13g2_a21o_1 _3484_ (.A2(_1904_),
    .A1(net984),
    .B1(_1878_),
    .X(_1905_));
 sg13g2_a21oi_1 _3485_ (.A1(net994),
    .A2(_1905_),
    .Y(_1906_),
    .B1(_1877_));
 sg13g2_nand2_1 _3486_ (.Y(_1907_),
    .A(net988),
    .B(net511));
 sg13g2_mux2_1 _3487_ (.A0(\s0.data_out[5][6] ),
    .A1(\s0.data_out[4][6] ),
    .S(net988),
    .X(_1908_));
 sg13g2_a21o_1 _3488_ (.A2(_1908_),
    .A1(net984),
    .B1(_1871_),
    .X(_1909_));
 sg13g2_a21oi_1 _3489_ (.A1(net996),
    .A2(_1909_),
    .Y(_1910_),
    .B1(_1870_));
 sg13g2_a22oi_1 _3490_ (.Y(_1911_),
    .B1(_1910_),
    .B2(net1240),
    .A2(_1906_),
    .A1(net1233));
 sg13g2_or2_1 _3491_ (.X(_1912_),
    .B(_1906_),
    .A(net1233));
 sg13g2_or2_1 _3492_ (.X(_1913_),
    .B(_1910_),
    .A(net1240));
 sg13g2_nand3_1 _3493_ (.B(_1912_),
    .C(_1913_),
    .A(_1911_),
    .Y(_1914_));
 sg13g2_mux2_1 _3494_ (.A0(\s0.data_out[5][4] ),
    .A1(\s0.data_out[4][4] ),
    .S(net989),
    .X(_1915_));
 sg13g2_a21oi_1 _3495_ (.A1(net982),
    .A2(_1915_),
    .Y(_1916_),
    .B1(_1858_));
 sg13g2_nand2b_1 _3496_ (.Y(_1917_),
    .B(net993),
    .A_N(_1916_));
 sg13g2_a21oi_1 _3497_ (.A1(_1856_),
    .A2(_1917_),
    .Y(_1918_),
    .B1(net1258));
 sg13g2_mux2_1 _3498_ (.A0(\s0.data_out[5][5] ),
    .A1(\s0.data_out[4][5] ),
    .S(net989),
    .X(_1919_));
 sg13g2_a21oi_1 _3499_ (.A1(net984),
    .A2(_1919_),
    .Y(_1920_),
    .B1(_1865_));
 sg13g2_nand2b_1 _3500_ (.Y(_1921_),
    .B(net994),
    .A_N(_1920_));
 sg13g2_nand3_1 _3501_ (.B(_1863_),
    .C(_1921_),
    .A(net1253),
    .Y(_1922_));
 sg13g2_nand2b_1 _3502_ (.Y(_1923_),
    .B(_1922_),
    .A_N(_1918_));
 sg13g2_a21oi_1 _3503_ (.A1(_1863_),
    .A2(_1921_),
    .Y(_1924_),
    .B1(net1253));
 sg13g2_nand3_1 _3504_ (.B(_1856_),
    .C(_1917_),
    .A(net1258),
    .Y(_1925_));
 sg13g2_o21ai_1 _3505_ (.B1(_1925_),
    .Y(_1926_),
    .A1(net1267),
    .A2(_1900_));
 sg13g2_nor4_1 _3506_ (.A(_1914_),
    .B(_1923_),
    .C(_1924_),
    .D(_1926_),
    .Y(_1927_));
 sg13g2_nand2_1 _3507_ (.Y(_1928_),
    .A(_1902_),
    .B(_1927_));
 sg13g2_o21ai_1 _3508_ (.B1(_1922_),
    .Y(_1929_),
    .A1(_1924_),
    .A2(_1925_));
 sg13g2_nor2b_1 _3509_ (.A(_1914_),
    .B_N(_1929_),
    .Y(_1930_));
 sg13g2_nor2b_1 _3510_ (.A(_1911_),
    .B_N(_1912_),
    .Y(_1931_));
 sg13g2_nor3_1 _3511_ (.A(_1821_),
    .B(_1930_),
    .C(_1931_),
    .Y(_1932_));
 sg13g2_or2_1 _3512_ (.X(_1933_),
    .B(net1208),
    .A(net318));
 sg13g2_a21oi_1 _3513_ (.A1(_1928_),
    .A2(_1932_),
    .Y(_0210_),
    .B1(_1933_));
 sg13g2_and2_1 _3514_ (.A(net1310),
    .B(net317),
    .X(_0211_));
 sg13g2_o21ai_1 _3515_ (.B1(net985),
    .Y(_1934_),
    .A1(net1226),
    .A2(net974));
 sg13g2_nand2_1 _3516_ (.Y(_1935_),
    .A(net1222),
    .B(net977));
 sg13g2_nand2b_1 _3517_ (.Y(_1936_),
    .B(_1935_),
    .A_N(_1934_));
 sg13g2_o21ai_1 _3518_ (.B1(_1936_),
    .Y(_1937_),
    .A1(net983),
    .A2(_1818_));
 sg13g2_nor2_1 _3519_ (.A(net353),
    .B(_1937_),
    .Y(_1938_));
 sg13g2_nor2_1 _3520_ (.A(net319),
    .B(net978),
    .Y(_1939_));
 sg13g2_nor2_1 _3521_ (.A(net972),
    .B(_1934_),
    .Y(_1940_));
 sg13g2_o21ai_1 _3522_ (.B1(_2471_),
    .Y(_1941_),
    .A1(net319),
    .A2(net988));
 sg13g2_o21ai_1 _3523_ (.B1(_1941_),
    .Y(_1942_),
    .A1(_1936_),
    .A2(_1939_));
 sg13g2_o21ai_1 _3524_ (.B1(net1313),
    .Y(_1943_),
    .A1(_1940_),
    .A2(_1942_));
 sg13g2_nor2_1 _3525_ (.A(_1938_),
    .B(_1943_),
    .Y(_0212_));
 sg13g2_nor2_1 _3526_ (.A(net1219),
    .B(_1937_),
    .Y(_0213_));
 sg13g2_mux2_1 _3527_ (.A0(\s0.data_out[3][0] ),
    .A1(\s0.data_out[4][0] ),
    .S(net987),
    .X(_1944_));
 sg13g2_nand2_1 _3528_ (.Y(_1945_),
    .A(net914),
    .B(_1944_));
 sg13g2_and2_1 _3529_ (.A(net969),
    .B(\s0.data_out[3][0] ),
    .X(_1946_));
 sg13g2_nor2b_1 _3530_ (.A(net969),
    .B_N(net1076),
    .Y(_1947_));
 sg13g2_o21ai_1 _3531_ (.B1(net980),
    .Y(_1948_),
    .A1(_1946_),
    .A2(_1947_));
 sg13g2_nand3_1 _3532_ (.B(_1945_),
    .C(_1948_),
    .A(net1308),
    .Y(_1949_));
 sg13g2_o21ai_1 _3533_ (.B1(_1949_),
    .Y(_1950_),
    .A1(net1308),
    .A2(net440));
 sg13g2_inv_1 _3534_ (.Y(_0214_),
    .A(_1950_));
 sg13g2_mux2_1 _3535_ (.A0(\s0.data_out[3][1] ),
    .A1(\s0.data_out[4][1] ),
    .S(net987),
    .X(_1951_));
 sg13g2_nand2_1 _3536_ (.Y(_1952_),
    .A(net914),
    .B(_1951_));
 sg13g2_and2_1 _3537_ (.A(net970),
    .B(\s0.data_out[3][1] ),
    .X(_1953_));
 sg13g2_nor2b_1 _3538_ (.A(net969),
    .B_N(net1072),
    .Y(_1954_));
 sg13g2_o21ai_1 _3539_ (.B1(net980),
    .Y(_1955_),
    .A1(_1953_),
    .A2(_1954_));
 sg13g2_nand3_1 _3540_ (.B(_1952_),
    .C(_1955_),
    .A(net1312),
    .Y(_1956_));
 sg13g2_o21ai_1 _3541_ (.B1(_1956_),
    .Y(_1957_),
    .A1(net1312),
    .A2(net433));
 sg13g2_inv_1 _3542_ (.Y(_0215_),
    .A(_1957_));
 sg13g2_nand2b_1 _3543_ (.Y(_1958_),
    .B(net420),
    .A_N(net987));
 sg13g2_a21oi_1 _3544_ (.A1(_1883_),
    .A2(_1958_),
    .Y(_1959_),
    .B1(net980));
 sg13g2_nor2b_1 _3545_ (.A(net969),
    .B_N(net1068),
    .Y(_1960_));
 sg13g2_a21oi_1 _3546_ (.A1(net969),
    .A2(net420),
    .Y(_1961_),
    .B1(_1960_));
 sg13g2_o21ai_1 _3547_ (.B1(net1312),
    .Y(_1962_),
    .A1(net914),
    .A2(_1961_));
 sg13g2_or2_1 _3548_ (.X(_1963_),
    .B(net533),
    .A(net1312));
 sg13g2_o21ai_1 _3549_ (.B1(_1963_),
    .Y(_1964_),
    .A1(_1959_),
    .A2(_1962_));
 sg13g2_inv_1 _3550_ (.Y(_0216_),
    .A(net534));
 sg13g2_mux2_1 _3551_ (.A0(\s0.data_out[3][3] ),
    .A1(\s0.data_out[4][3] ),
    .S(net987),
    .X(_1965_));
 sg13g2_nand2_1 _3552_ (.Y(_1966_),
    .A(net914),
    .B(_1965_));
 sg13g2_and2_1 _3553_ (.A(net970),
    .B(\s0.data_out[3][3] ),
    .X(_1967_));
 sg13g2_nor2b_1 _3554_ (.A(net970),
    .B_N(net1064),
    .Y(_1968_));
 sg13g2_o21ai_1 _3555_ (.B1(net980),
    .Y(_1969_),
    .A1(_1967_),
    .A2(_1968_));
 sg13g2_nand3_1 _3556_ (.B(_1966_),
    .C(_1969_),
    .A(net1312),
    .Y(_1970_));
 sg13g2_o21ai_1 _3557_ (.B1(_1970_),
    .Y(_1971_),
    .A1(net1312),
    .A2(net403));
 sg13g2_inv_1 _3558_ (.Y(_0217_),
    .A(_1971_));
 sg13g2_mux2_1 _3559_ (.A0(\s0.data_out[3][4] ),
    .A1(\s0.data_out[4][4] ),
    .S(net987),
    .X(_1972_));
 sg13g2_nand2_1 _3560_ (.Y(_1973_),
    .A(net914),
    .B(_1972_));
 sg13g2_and2_1 _3561_ (.A(net970),
    .B(\s0.data_out[3][4] ),
    .X(_1974_));
 sg13g2_nor2b_1 _3562_ (.A(net970),
    .B_N(net1058),
    .Y(_1975_));
 sg13g2_o21ai_1 _3563_ (.B1(net986),
    .Y(_1976_),
    .A1(_1974_),
    .A2(_1975_));
 sg13g2_nand3_1 _3564_ (.B(_1973_),
    .C(_1976_),
    .A(net1308),
    .Y(_1977_));
 sg13g2_o21ai_1 _3565_ (.B1(_1977_),
    .Y(_1978_),
    .A1(net1308),
    .A2(net443));
 sg13g2_inv_1 _3566_ (.Y(_0218_),
    .A(net444));
 sg13g2_mux2_1 _3567_ (.A0(\s0.data_out[3][5] ),
    .A1(\s0.data_out[4][5] ),
    .S(net988),
    .X(_1979_));
 sg13g2_nand2_1 _3568_ (.Y(_1980_),
    .A(_2471_),
    .B(_1979_));
 sg13g2_and2_1 _3569_ (.A(net972),
    .B(\s0.data_out[3][5] ),
    .X(_1981_));
 sg13g2_nor2b_1 _3570_ (.A(net972),
    .B_N(net1054),
    .Y(_1982_));
 sg13g2_o21ai_1 _3571_ (.B1(net983),
    .Y(_1983_),
    .A1(_1981_),
    .A2(_1982_));
 sg13g2_nand3_1 _3572_ (.B(_1980_),
    .C(_1983_),
    .A(net1313),
    .Y(_1984_));
 sg13g2_o21ai_1 _3573_ (.B1(_1984_),
    .Y(_1985_),
    .A1(net1313),
    .A2(net470));
 sg13g2_inv_1 _3574_ (.Y(_0219_),
    .A(_1985_));
 sg13g2_nand2b_1 _3575_ (.Y(_1986_),
    .B(\s0.data_out[3][6] ),
    .A_N(net988));
 sg13g2_a21oi_1 _3576_ (.A1(_1907_),
    .A2(_1986_),
    .Y(_1987_),
    .B1(net983));
 sg13g2_nor2b_1 _3577_ (.A(net974),
    .B_N(net1050),
    .Y(_1988_));
 sg13g2_a21oi_1 _3578_ (.A1(net972),
    .A2(\s0.data_out[3][6] ),
    .Y(_1989_),
    .B1(_1988_));
 sg13g2_o21ai_1 _3579_ (.B1(net1310),
    .Y(_1990_),
    .A1(net914),
    .A2(_1989_));
 sg13g2_or2_1 _3580_ (.X(_1991_),
    .B(net511),
    .A(net1313));
 sg13g2_o21ai_1 _3581_ (.B1(_1991_),
    .Y(_1992_),
    .A1(_1987_),
    .A2(_1990_));
 sg13g2_inv_1 _3582_ (.Y(_0220_),
    .A(net512));
 sg13g2_nand2b_1 _3583_ (.Y(_1993_),
    .B(net515),
    .A_N(net988));
 sg13g2_a21oi_1 _3584_ (.A1(_1903_),
    .A2(_1993_),
    .Y(_1994_),
    .B1(net983));
 sg13g2_nor2b_1 _3585_ (.A(net974),
    .B_N(net1046),
    .Y(_1995_));
 sg13g2_a21oi_1 _3586_ (.A1(net972),
    .A2(net515),
    .Y(_1996_),
    .B1(_1995_));
 sg13g2_o21ai_1 _3587_ (.B1(net1309),
    .Y(_1997_),
    .A1(net914),
    .A2(_1996_));
 sg13g2_or2_1 _3588_ (.X(_1998_),
    .B(net535),
    .A(net1313));
 sg13g2_o21ai_1 _3589_ (.B1(_1998_),
    .Y(_1999_),
    .A1(_1994_),
    .A2(_1997_));
 sg13g2_inv_1 _3590_ (.Y(_0221_),
    .A(_1999_));
 sg13g2_mux2_1 _3591_ (.A0(\s0.data_out[4][2] ),
    .A1(\s0.data_out[3][2] ),
    .S(net979),
    .X(_2000_));
 sg13g2_a21o_1 _3592_ (.A2(_2000_),
    .A1(net969),
    .B1(_1960_),
    .X(_2001_));
 sg13g2_a21oi_1 _3593_ (.A1(net980),
    .A2(_2001_),
    .Y(_2002_),
    .B1(_1959_));
 sg13g2_or2_1 _3594_ (.X(_2003_),
    .B(_2002_),
    .A(net1269));
 sg13g2_mux2_1 _3595_ (.A0(\s0.data_out[4][1] ),
    .A1(\s0.data_out[3][1] ),
    .S(net976),
    .X(_2004_));
 sg13g2_a21oi_1 _3596_ (.A1(net969),
    .A2(_2004_),
    .Y(_2005_),
    .B1(_1954_));
 sg13g2_nand2b_1 _3597_ (.Y(_2006_),
    .B(net980),
    .A_N(_2005_));
 sg13g2_and2_1 _3598_ (.A(_1952_),
    .B(_2006_),
    .X(_2007_));
 sg13g2_mux2_1 _3599_ (.A0(\s0.data_out[4][0] ),
    .A1(\s0.data_out[3][0] ),
    .S(net976),
    .X(_2008_));
 sg13g2_a21oi_1 _3600_ (.A1(net969),
    .A2(_2008_),
    .Y(_2009_),
    .B1(_1947_));
 sg13g2_nand2b_1 _3601_ (.Y(_2010_),
    .B(net980),
    .A_N(_2009_));
 sg13g2_o21ai_1 _3602_ (.B1(_2003_),
    .Y(_2011_),
    .A1(net1275),
    .A2(_2007_));
 sg13g2_a221oi_1 _3603_ (.B2(_1945_),
    .C1(net1284),
    .B1(_2010_),
    .A1(net1275),
    .Y(_2012_),
    .A2(_2007_));
 sg13g2_nand2_1 _3604_ (.Y(_2013_),
    .A(net976),
    .B(net509));
 sg13g2_mux2_1 _3605_ (.A0(\s0.data_out[4][3] ),
    .A1(\s0.data_out[3][3] ),
    .S(net979),
    .X(_2014_));
 sg13g2_a21oi_1 _3606_ (.A1(net970),
    .A2(_2014_),
    .Y(_2015_),
    .B1(_1968_));
 sg13g2_nand2b_1 _3607_ (.Y(_2016_),
    .B(net980),
    .A_N(_2015_));
 sg13g2_and2_1 _3608_ (.A(_1966_),
    .B(_2016_),
    .X(_2017_));
 sg13g2_a22oi_1 _3609_ (.Y(_2018_),
    .B1(_2017_),
    .B2(net1263),
    .A2(_2002_),
    .A1(net1269));
 sg13g2_o21ai_1 _3610_ (.B1(_2018_),
    .Y(_2019_),
    .A1(_2011_),
    .A2(_2012_));
 sg13g2_nand2_1 _3611_ (.Y(_2020_),
    .A(net977),
    .B(net515));
 sg13g2_mux2_1 _3612_ (.A0(\s0.data_out[4][7] ),
    .A1(\s0.data_out[3][7] ),
    .S(net978),
    .X(_2021_));
 sg13g2_a21o_1 _3613_ (.A2(_2021_),
    .A1(net972),
    .B1(_1995_),
    .X(_2022_));
 sg13g2_a21oi_1 _3614_ (.A1(net983),
    .A2(_2022_),
    .Y(_2023_),
    .B1(_1994_));
 sg13g2_nand2_1 _3615_ (.Y(_2024_),
    .A(net977),
    .B(net576));
 sg13g2_mux2_1 _3616_ (.A0(\s0.data_out[4][6] ),
    .A1(\s0.data_out[3][6] ),
    .S(net978),
    .X(_2025_));
 sg13g2_a21o_1 _3617_ (.A2(_2025_),
    .A1(net972),
    .B1(_1988_),
    .X(_2026_));
 sg13g2_a21oi_1 _3618_ (.A1(net983),
    .A2(_2026_),
    .Y(_2027_),
    .B1(_1987_));
 sg13g2_a22oi_1 _3619_ (.Y(_2028_),
    .B1(_2027_),
    .B2(net1241),
    .A2(_2023_),
    .A1(net1233));
 sg13g2_or2_1 _3620_ (.X(_2029_),
    .B(_2027_),
    .A(net1241));
 sg13g2_or2_1 _3621_ (.X(_2030_),
    .B(_2023_),
    .A(net1234));
 sg13g2_and3_1 _3622_ (.X(_2031_),
    .A(_2028_),
    .B(_2029_),
    .C(_2030_));
 sg13g2_nand2_1 _3623_ (.Y(_2032_),
    .A(net977),
    .B(net355));
 sg13g2_mux2_1 _3624_ (.A0(\s0.data_out[4][5] ),
    .A1(\s0.data_out[3][5] ),
    .S(net978),
    .X(_2033_));
 sg13g2_a21oi_1 _3625_ (.A1(net972),
    .A2(_2033_),
    .Y(_2034_),
    .B1(_1982_));
 sg13g2_nand2b_1 _3626_ (.Y(_2035_),
    .B(net983),
    .A_N(_2034_));
 sg13g2_nand3_1 _3627_ (.B(_1980_),
    .C(_2035_),
    .A(net1249),
    .Y(_2036_));
 sg13g2_o21ai_1 _3628_ (.B1(_2036_),
    .Y(_2037_),
    .A1(net1263),
    .A2(_2017_));
 sg13g2_mux2_1 _3629_ (.A0(\s0.data_out[4][4] ),
    .A1(\s0.data_out[3][4] ),
    .S(net979),
    .X(_2038_));
 sg13g2_a21oi_1 _3630_ (.A1(net970),
    .A2(_2038_),
    .Y(_2039_),
    .B1(_1975_));
 sg13g2_o21ai_1 _3631_ (.B1(_1973_),
    .Y(_2040_),
    .A1(net914),
    .A2(_2039_));
 sg13g2_or2_1 _3632_ (.X(_2041_),
    .B(_2040_),
    .A(net1215));
 sg13g2_xnor2_1 _3633_ (.Y(_2042_),
    .A(net1215),
    .B(_2040_));
 sg13g2_a21oi_1 _3634_ (.A1(_1980_),
    .A2(_2035_),
    .Y(_2043_),
    .B1(net1249));
 sg13g2_nor3_1 _3635_ (.A(_2037_),
    .B(_2042_),
    .C(_2043_),
    .Y(_2044_));
 sg13g2_nand3_1 _3636_ (.B(_2031_),
    .C(_2044_),
    .A(_2019_),
    .Y(_2045_));
 sg13g2_o21ai_1 _3637_ (.B1(_2036_),
    .Y(_2046_),
    .A1(_2041_),
    .A2(_2043_));
 sg13g2_nand2b_1 _3638_ (.Y(_2047_),
    .B(_2030_),
    .A_N(_2028_));
 sg13g2_a21oi_1 _3639_ (.A1(_2031_),
    .A2(_2046_),
    .Y(_2048_),
    .B1(_1937_));
 sg13g2_and2_1 _3640_ (.A(_2047_),
    .B(_2048_),
    .X(_2049_));
 sg13g2_or2_1 _3641_ (.X(_2050_),
    .B(net1210),
    .A(net317));
 sg13g2_a21oi_1 _3642_ (.A1(_2045_),
    .A2(_2049_),
    .Y(_0222_),
    .B1(_2050_));
 sg13g2_and2_1 _3643_ (.A(net1309),
    .B(net311),
    .X(_0223_));
 sg13g2_o21ai_1 _3644_ (.B1(net973),
    .Y(_2051_),
    .A1(net1227),
    .A2(net963));
 sg13g2_nor2b_1 _3645_ (.A(net1227),
    .B_N(net967),
    .Y(_2052_));
 sg13g2_nor2_1 _3646_ (.A(_2051_),
    .B(_2052_),
    .Y(_2053_));
 sg13g2_a21oi_1 _3647_ (.A1(net932),
    .A2(_1935_),
    .Y(_2054_),
    .B1(_2053_));
 sg13g2_inv_1 _3648_ (.Y(_2055_),
    .A(_2054_));
 sg13g2_o21ai_1 _3649_ (.B1(_2053_),
    .Y(_2056_),
    .A1(\s0.was_valid_out[2] [0]),
    .A2(net967));
 sg13g2_nor2_1 _3650_ (.A(net963),
    .B(_2051_),
    .Y(_2057_));
 sg13g2_o21ai_1 _3651_ (.B1(net933),
    .Y(_2058_),
    .A1(\s0.was_valid_out[2] [0]),
    .A2(net977));
 sg13g2_nand2_1 _3652_ (.Y(_2059_),
    .A(_2056_),
    .B(_2058_));
 sg13g2_o21ai_1 _3653_ (.B1(net1309),
    .Y(_2060_),
    .A1(_2057_),
    .A2(_2059_));
 sg13g2_a21oi_1 _3654_ (.A1(_2443_),
    .A2(_2054_),
    .Y(_0224_),
    .B1(_2060_));
 sg13g2_nor2_1 _3655_ (.A(net1219),
    .B(_2055_),
    .Y(_0225_));
 sg13g2_mux2_1 _3656_ (.A0(\s0.data_out[2][0] ),
    .A1(\s0.data_out[3][0] ),
    .S(net976),
    .X(_2061_));
 sg13g2_nand2_1 _3657_ (.Y(_2062_),
    .A(net932),
    .B(_2061_));
 sg13g2_and2_1 _3658_ (.A(net959),
    .B(\s0.data_out[2][0] ),
    .X(_2063_));
 sg13g2_nor2b_1 _3659_ (.A(net959),
    .B_N(net1076),
    .Y(_2064_));
 sg13g2_o21ai_1 _3660_ (.B1(net971),
    .Y(_2065_),
    .A1(_2063_),
    .A2(_2064_));
 sg13g2_nand3_1 _3661_ (.B(_2062_),
    .C(_2065_),
    .A(net1307),
    .Y(_2066_));
 sg13g2_o21ai_1 _3662_ (.B1(_2066_),
    .Y(_2067_),
    .A1(net1297),
    .A2(net437));
 sg13g2_inv_1 _3663_ (.Y(_0226_),
    .A(_2067_));
 sg13g2_mux2_1 _3664_ (.A0(\s0.data_out[2][1] ),
    .A1(\s0.data_out[3][1] ),
    .S(net976),
    .X(_2068_));
 sg13g2_nand2_1 _3665_ (.Y(_2069_),
    .A(net932),
    .B(_2068_));
 sg13g2_and2_1 _3666_ (.A(net960),
    .B(\s0.data_out[2][1] ),
    .X(_2070_));
 sg13g2_nor2b_1 _3667_ (.A(net959),
    .B_N(net1072),
    .Y(_2071_));
 sg13g2_o21ai_1 _3668_ (.B1(net971),
    .Y(_2072_),
    .A1(_2070_),
    .A2(_2071_));
 sg13g2_nand3_1 _3669_ (.B(_2069_),
    .C(_2072_),
    .A(net1307),
    .Y(_2073_));
 sg13g2_o21ai_1 _3670_ (.B1(_2073_),
    .Y(_2074_),
    .A1(net1307),
    .A2(net421));
 sg13g2_inv_1 _3671_ (.Y(_0227_),
    .A(_2074_));
 sg13g2_mux2_1 _3672_ (.A0(\s0.data_out[2][2] ),
    .A1(\s0.data_out[3][2] ),
    .S(net976),
    .X(_2075_));
 sg13g2_nand2_1 _3673_ (.Y(_2076_),
    .A(net932),
    .B(_2075_));
 sg13g2_and2_1 _3674_ (.A(net959),
    .B(net611),
    .X(_2077_));
 sg13g2_nor2b_1 _3675_ (.A(net959),
    .B_N(net1068),
    .Y(_2078_));
 sg13g2_o21ai_1 _3676_ (.B1(net971),
    .Y(_2079_),
    .A1(_2077_),
    .A2(_2078_));
 sg13g2_nand3_1 _3677_ (.B(_2076_),
    .C(_2079_),
    .A(net1307),
    .Y(_2080_));
 sg13g2_o21ai_1 _3678_ (.B1(_2080_),
    .Y(_2081_),
    .A1(net1307),
    .A2(net420));
 sg13g2_inv_1 _3679_ (.Y(_0228_),
    .A(_2081_));
 sg13g2_nand2b_1 _3680_ (.Y(_2082_),
    .B(net446),
    .A_N(net976));
 sg13g2_a21oi_1 _3681_ (.A1(_2013_),
    .A2(_2082_),
    .Y(_2083_),
    .B1(net971));
 sg13g2_nor2b_1 _3682_ (.A(net960),
    .B_N(net1064),
    .Y(_2084_));
 sg13g2_a21oi_1 _3683_ (.A1(net960),
    .A2(net446),
    .Y(_2085_),
    .B1(_2084_));
 sg13g2_o21ai_1 _3684_ (.B1(net1307),
    .Y(_2086_),
    .A1(net932),
    .A2(_2085_));
 sg13g2_or2_1 _3685_ (.X(_2087_),
    .B(net509),
    .A(net1308));
 sg13g2_o21ai_1 _3686_ (.B1(_2087_),
    .Y(_2088_),
    .A1(_2083_),
    .A2(_2086_));
 sg13g2_inv_1 _3687_ (.Y(_0229_),
    .A(net510));
 sg13g2_mux2_1 _3688_ (.A0(\s0.data_out[2][4] ),
    .A1(\s0.data_out[3][4] ),
    .S(net976),
    .X(_2089_));
 sg13g2_nand2_1 _3689_ (.Y(_2090_),
    .A(net932),
    .B(_2089_));
 sg13g2_and2_1 _3690_ (.A(net960),
    .B(\s0.data_out[2][4] ),
    .X(_2091_));
 sg13g2_nor2b_1 _3691_ (.A(net960),
    .B_N(net1058),
    .Y(_2092_));
 sg13g2_o21ai_1 _3692_ (.B1(net971),
    .Y(_2093_),
    .A1(_2091_),
    .A2(_2092_));
 sg13g2_nand3_1 _3693_ (.B(_2090_),
    .C(_2093_),
    .A(net1307),
    .Y(_2094_));
 sg13g2_o21ai_1 _3694_ (.B1(_2094_),
    .Y(_2095_),
    .A1(net1307),
    .A2(net441));
 sg13g2_inv_1 _3695_ (.Y(_0230_),
    .A(_2095_));
 sg13g2_nand2b_1 _3696_ (.Y(_2096_),
    .B(net349),
    .A_N(net977));
 sg13g2_a21oi_1 _3697_ (.A1(_2032_),
    .A2(_2096_),
    .Y(_2097_),
    .B1(net973));
 sg13g2_nor2b_1 _3698_ (.A(net963),
    .B_N(net1054),
    .Y(_2098_));
 sg13g2_a21oi_1 _3699_ (.A1(net963),
    .A2(net349),
    .Y(_2099_),
    .B1(_2098_));
 sg13g2_o21ai_1 _3700_ (.B1(net1309),
    .Y(_2100_),
    .A1(net933),
    .A2(_2099_));
 sg13g2_or2_1 _3701_ (.X(_2101_),
    .B(net355),
    .A(net1310));
 sg13g2_o21ai_1 _3702_ (.B1(_2101_),
    .Y(_2102_),
    .A1(_2097_),
    .A2(_2100_));
 sg13g2_inv_1 _3703_ (.Y(_0231_),
    .A(_2102_));
 sg13g2_nand2b_1 _3704_ (.Y(_2103_),
    .B(net491),
    .A_N(net977));
 sg13g2_a21oi_1 _3705_ (.A1(_2024_),
    .A2(_2103_),
    .Y(_2104_),
    .B1(net973));
 sg13g2_nor2b_1 _3706_ (.A(net964),
    .B_N(net1050),
    .Y(_2105_));
 sg13g2_a21oi_1 _3707_ (.A1(net964),
    .A2(net491),
    .Y(_2106_),
    .B1(_2105_));
 sg13g2_o21ai_1 _3708_ (.B1(net1309),
    .Y(_2107_),
    .A1(net933),
    .A2(_2106_));
 sg13g2_or2_1 _3709_ (.X(_2108_),
    .B(net576),
    .A(net1309));
 sg13g2_o21ai_1 _3710_ (.B1(_2108_),
    .Y(_2109_),
    .A1(_2104_),
    .A2(_2107_));
 sg13g2_inv_1 _3711_ (.Y(_0232_),
    .A(_2109_));
 sg13g2_nand2b_1 _3712_ (.Y(_2110_),
    .B(\s0.data_out[2][7] ),
    .A_N(net977));
 sg13g2_a21oi_1 _3713_ (.A1(_2020_),
    .A2(_2110_),
    .Y(_2111_),
    .B1(net973));
 sg13g2_nor2b_1 _3714_ (.A(net963),
    .B_N(net1046),
    .Y(_2112_));
 sg13g2_a21oi_1 _3715_ (.A1(net963),
    .A2(\s0.data_out[2][7] ),
    .Y(_2113_),
    .B1(_2112_));
 sg13g2_o21ai_1 _3716_ (.B1(net1309),
    .Y(_2114_),
    .A1(net933),
    .A2(_2113_));
 sg13g2_or2_1 _3717_ (.X(_2115_),
    .B(net515),
    .A(net1309));
 sg13g2_o21ai_1 _3718_ (.B1(_2115_),
    .Y(_2116_),
    .A1(_2111_),
    .A2(_2114_));
 sg13g2_inv_1 _3719_ (.Y(_0233_),
    .A(net516));
 sg13g2_nand2_1 _3720_ (.Y(_2117_),
    .A(net968),
    .B(net488));
 sg13g2_o21ai_1 _3721_ (.B1(_2117_),
    .Y(_2118_),
    .A1(net968),
    .A2(_2492_));
 sg13g2_a21oi_1 _3722_ (.A1(net959),
    .A2(_2118_),
    .Y(_2119_),
    .B1(_2078_));
 sg13g2_o21ai_1 _3723_ (.B1(_2076_),
    .Y(_2120_),
    .A1(net932),
    .A2(_2119_));
 sg13g2_mux2_1 _3724_ (.A0(\s0.data_out[3][1] ),
    .A1(\s0.data_out[2][1] ),
    .S(net965),
    .X(_2121_));
 sg13g2_a21oi_1 _3725_ (.A1(net959),
    .A2(_2121_),
    .Y(_2122_),
    .B1(_2071_));
 sg13g2_nand2b_1 _3726_ (.Y(_2123_),
    .B(net971),
    .A_N(_2122_));
 sg13g2_nand3_1 _3727_ (.B(_2069_),
    .C(_2123_),
    .A(net1275),
    .Y(_2124_));
 sg13g2_mux2_1 _3728_ (.A0(\s0.data_out[3][0] ),
    .A1(\s0.data_out[2][0] ),
    .S(net965),
    .X(_2125_));
 sg13g2_a21oi_1 _3729_ (.A1(net959),
    .A2(_2125_),
    .Y(_2126_),
    .B1(_2064_));
 sg13g2_o21ai_1 _3730_ (.B1(_2062_),
    .Y(_2127_),
    .A1(net932),
    .A2(_2126_));
 sg13g2_nor2b_1 _3731_ (.A(net1284),
    .B_N(_2127_),
    .Y(_2128_));
 sg13g2_a21oi_1 _3732_ (.A1(_2069_),
    .A2(_2123_),
    .Y(_2129_),
    .B1(net1276));
 sg13g2_a221oi_1 _3733_ (.B2(_2128_),
    .C1(_2129_),
    .B1(_2124_),
    .A1(net1212),
    .Y(_2130_),
    .A2(_2120_));
 sg13g2_mux2_1 _3734_ (.A0(\s0.data_out[3][3] ),
    .A1(\s0.data_out[2][3] ),
    .S(net965),
    .X(_2131_));
 sg13g2_a21o_1 _3735_ (.A2(_2131_),
    .A1(net960),
    .B1(_2084_),
    .X(_2132_));
 sg13g2_a21oi_1 _3736_ (.A1(net971),
    .A2(_2132_),
    .Y(_2133_),
    .B1(_2083_));
 sg13g2_nand2_1 _3737_ (.Y(_2134_),
    .A(net1262),
    .B(_2133_));
 sg13g2_o21ai_1 _3738_ (.B1(_2134_),
    .Y(_2135_),
    .A1(net1211),
    .A2(_2120_));
 sg13g2_nand2_1 _3739_ (.Y(_2136_),
    .A(net966),
    .B(net553));
 sg13g2_mux2_1 _3740_ (.A0(\s0.data_out[3][7] ),
    .A1(\s0.data_out[2][7] ),
    .S(net967),
    .X(_2137_));
 sg13g2_a21o_1 _3741_ (.A2(_2137_),
    .A1(net963),
    .B1(_2112_),
    .X(_2138_));
 sg13g2_a21oi_1 _3742_ (.A1(net973),
    .A2(_2138_),
    .Y(_2139_),
    .B1(_2111_));
 sg13g2_nand2_1 _3743_ (.Y(_2140_),
    .A(net966),
    .B(net491));
 sg13g2_mux2_1 _3744_ (.A0(\s0.data_out[3][6] ),
    .A1(\s0.data_out[2][6] ),
    .S(net967),
    .X(_2141_));
 sg13g2_a21o_1 _3745_ (.A2(_2141_),
    .A1(net964),
    .B1(_2105_),
    .X(_2142_));
 sg13g2_a21oi_1 _3746_ (.A1(net973),
    .A2(_2142_),
    .Y(_2143_),
    .B1(_2104_));
 sg13g2_a22oi_1 _3747_ (.Y(_2144_),
    .B1(_2143_),
    .B2(net1240),
    .A2(_2139_),
    .A1(net1233));
 sg13g2_nor2_1 _3748_ (.A(net1241),
    .B(_2143_),
    .Y(_2145_));
 sg13g2_or2_1 _3749_ (.X(_2146_),
    .B(_2139_),
    .A(net1234));
 sg13g2_nand3b_1 _3750_ (.B(_2146_),
    .C(_2144_),
    .Y(_2147_),
    .A_N(_2145_));
 sg13g2_mux2_1 _3751_ (.A0(\s0.data_out[3][4] ),
    .A1(\s0.data_out[2][4] ),
    .S(net965),
    .X(_2148_));
 sg13g2_a21oi_1 _3752_ (.A1(net960),
    .A2(_2148_),
    .Y(_2149_),
    .B1(_2092_));
 sg13g2_nand2b_1 _3753_ (.Y(_2150_),
    .B(net971),
    .A_N(_2149_));
 sg13g2_and2_1 _3754_ (.A(_2090_),
    .B(_2150_),
    .X(_2151_));
 sg13g2_mux2_1 _3755_ (.A0(\s0.data_out[3][5] ),
    .A1(\s0.data_out[2][5] ),
    .S(net966),
    .X(_2152_));
 sg13g2_a21o_1 _3756_ (.A2(_2152_),
    .A1(net963),
    .B1(_2098_),
    .X(_2153_));
 sg13g2_a21oi_1 _3757_ (.A1(net973),
    .A2(_2153_),
    .Y(_2154_),
    .B1(_2097_));
 sg13g2_a22oi_1 _3758_ (.Y(_2155_),
    .B1(_2154_),
    .B2(net1248),
    .A2(_2151_),
    .A1(net1255));
 sg13g2_nor2_1 _3759_ (.A(net1248),
    .B(_2154_),
    .Y(_2156_));
 sg13g2_nor2_1 _3760_ (.A(net1262),
    .B(_2133_),
    .Y(_2157_));
 sg13g2_nor2_1 _3761_ (.A(_2156_),
    .B(_2157_),
    .Y(_2158_));
 sg13g2_o21ai_1 _3762_ (.B1(_2155_),
    .Y(_2159_),
    .A1(net1255),
    .A2(_2151_));
 sg13g2_o21ai_1 _3763_ (.B1(_2158_),
    .Y(_2160_),
    .A1(_2130_),
    .A2(_2135_));
 sg13g2_or3_1 _3764_ (.A(_2147_),
    .B(_2159_),
    .C(_2160_),
    .X(_2161_));
 sg13g2_nor3_1 _3765_ (.A(_2147_),
    .B(_2155_),
    .C(_2156_),
    .Y(_2162_));
 sg13g2_nor2b_1 _3766_ (.A(_2144_),
    .B_N(_2146_),
    .Y(_2163_));
 sg13g2_nor3_1 _3767_ (.A(_2055_),
    .B(_2162_),
    .C(_2163_),
    .Y(_2164_));
 sg13g2_or2_1 _3768_ (.X(_2165_),
    .B(net1210),
    .A(net311));
 sg13g2_a21oi_1 _3769_ (.A1(_2161_),
    .A2(_2164_),
    .Y(_0234_),
    .B1(_2165_));
 sg13g2_and2_1 _3770_ (.A(net1298),
    .B(net300),
    .X(_0235_));
 sg13g2_o21ai_1 _3771_ (.B1(net962),
    .Y(_2166_),
    .A1(net1225),
    .A2(net953));
 sg13g2_nand2_1 _3772_ (.Y(_2167_),
    .A(net1222),
    .B(net956));
 sg13g2_a21oi_1 _3773_ (.A1(net1222),
    .A2(net957),
    .Y(_2168_),
    .B1(_2166_));
 sg13g2_inv_1 _3774_ (.Y(_2169_),
    .A(_2168_));
 sg13g2_o21ai_1 _3775_ (.B1(_2169_),
    .Y(_2170_),
    .A1(net962),
    .A2(_2052_));
 sg13g2_o21ai_1 _3776_ (.B1(_2168_),
    .Y(_2171_),
    .A1(net328),
    .A2(net957));
 sg13g2_o21ai_1 _3777_ (.B1(net930),
    .Y(_2172_),
    .A1(net328),
    .A2(net966));
 sg13g2_o21ai_1 _3778_ (.B1(_2172_),
    .Y(_2173_),
    .A1(net953),
    .A2(_2166_));
 sg13g2_inv_1 _3779_ (.Y(_2174_),
    .A(_2173_));
 sg13g2_o21ai_1 _3780_ (.B1(net1299),
    .Y(_2175_),
    .A1(net393),
    .A2(_2170_));
 sg13g2_a21oi_1 _3781_ (.A1(_2171_),
    .A2(_2174_),
    .Y(_0236_),
    .B1(_2175_));
 sg13g2_nor2_1 _3782_ (.A(net1218),
    .B(_2170_),
    .Y(_0237_));
 sg13g2_mux2_1 _3783_ (.A0(\s0.data_out[1][0] ),
    .A1(\s0.data_out[2][0] ),
    .S(net965),
    .X(_2176_));
 sg13g2_nand2_1 _3784_ (.Y(_2177_),
    .A(net930),
    .B(_2176_));
 sg13g2_and2_1 _3785_ (.A(net949),
    .B(\s0.data_out[1][0] ),
    .X(_2178_));
 sg13g2_nor2b_1 _3786_ (.A(net949),
    .B_N(net1073),
    .Y(_2179_));
 sg13g2_o21ai_1 _3787_ (.B1(net961),
    .Y(_2180_),
    .A1(_2178_),
    .A2(_2179_));
 sg13g2_nand3_1 _3788_ (.B(_2177_),
    .C(_2180_),
    .A(net1297),
    .Y(_2181_));
 sg13g2_o21ai_1 _3789_ (.B1(_2181_),
    .Y(_2182_),
    .A1(net1300),
    .A2(net424));
 sg13g2_inv_1 _3790_ (.Y(_0238_),
    .A(net425));
 sg13g2_mux2_1 _3791_ (.A0(\s0.data_out[1][1] ),
    .A1(\s0.data_out[2][1] ),
    .S(net965),
    .X(_2183_));
 sg13g2_nand2_1 _3792_ (.Y(_2184_),
    .A(net930),
    .B(_2183_));
 sg13g2_and2_1 _3793_ (.A(net949),
    .B(\s0.data_out[1][1] ),
    .X(_2185_));
 sg13g2_nor2b_1 _3794_ (.A(net949),
    .B_N(net1069),
    .Y(_2186_));
 sg13g2_o21ai_1 _3795_ (.B1(net961),
    .Y(_2187_),
    .A1(_2185_),
    .A2(_2186_));
 sg13g2_nand3_1 _3796_ (.B(_2184_),
    .C(_2187_),
    .A(net1297),
    .Y(_2188_));
 sg13g2_o21ai_1 _3797_ (.B1(_2188_),
    .Y(_2189_),
    .A1(net1297),
    .A2(net426));
 sg13g2_inv_1 _3798_ (.Y(_0239_),
    .A(net427));
 sg13g2_nand2b_1 _3799_ (.Y(_2190_),
    .B(net458),
    .A_N(net965));
 sg13g2_a21oi_1 _3800_ (.A1(_2117_),
    .A2(_2190_),
    .Y(_2191_),
    .B1(net961));
 sg13g2_nor2b_1 _3801_ (.A(net949),
    .B_N(net1065),
    .Y(_2192_));
 sg13g2_a21oi_1 _3802_ (.A1(net949),
    .A2(net458),
    .Y(_2193_),
    .B1(_2192_));
 sg13g2_o21ai_1 _3803_ (.B1(net1297),
    .Y(_2194_),
    .A1(net930),
    .A2(_2193_));
 sg13g2_or2_1 _3804_ (.X(_2195_),
    .B(net488),
    .A(net1297));
 sg13g2_o21ai_1 _3805_ (.B1(_2195_),
    .Y(_2196_),
    .A1(_2191_),
    .A2(_2194_));
 sg13g2_inv_1 _3806_ (.Y(_0240_),
    .A(net489));
 sg13g2_mux2_1 _3807_ (.A0(\s0.data_out[1][3] ),
    .A1(\s0.data_out[2][3] ),
    .S(net965),
    .X(_2197_));
 sg13g2_nand2_1 _3808_ (.Y(_2198_),
    .A(net930),
    .B(_2197_));
 sg13g2_and2_1 _3809_ (.A(net950),
    .B(\s0.data_out[1][3] ),
    .X(_2199_));
 sg13g2_nor2b_1 _3810_ (.A(net950),
    .B_N(net1061),
    .Y(_2200_));
 sg13g2_o21ai_1 _3811_ (.B1(net961),
    .Y(_2201_),
    .A1(_2199_),
    .A2(_2200_));
 sg13g2_nand3_1 _3812_ (.B(_2198_),
    .C(_2201_),
    .A(net1297),
    .Y(_2202_));
 sg13g2_o21ai_1 _3813_ (.B1(_2202_),
    .Y(_2203_),
    .A1(net1297),
    .A2(net446));
 sg13g2_inv_1 _3814_ (.Y(_0241_),
    .A(net447));
 sg13g2_mux2_1 _3815_ (.A0(\s0.data_out[1][4] ),
    .A1(\s0.data_out[2][4] ),
    .S(net966),
    .X(_2204_));
 sg13g2_nand2_1 _3816_ (.Y(_2205_),
    .A(net930),
    .B(_2204_));
 sg13g2_and2_1 _3817_ (.A(net950),
    .B(\s0.data_out[1][4] ),
    .X(_2206_));
 sg13g2_nor2b_1 _3818_ (.A(net950),
    .B_N(net1057),
    .Y(_2207_));
 sg13g2_o21ai_1 _3819_ (.B1(net962),
    .Y(_2208_),
    .A1(_2206_),
    .A2(_2207_));
 sg13g2_nand3_1 _3820_ (.B(_2205_),
    .C(_2208_),
    .A(net1298),
    .Y(_2209_));
 sg13g2_o21ai_1 _3821_ (.B1(_2209_),
    .Y(_2210_),
    .A1(net1298),
    .A2(net417));
 sg13g2_inv_1 _3822_ (.Y(_0242_),
    .A(_2210_));
 sg13g2_mux2_1 _3823_ (.A0(\s0.data_out[1][5] ),
    .A1(\s0.data_out[2][5] ),
    .S(net966),
    .X(_2211_));
 sg13g2_nand2_1 _3824_ (.Y(_2212_),
    .A(net930),
    .B(_2211_));
 sg13g2_and2_1 _3825_ (.A(net953),
    .B(\s0.data_out[1][5] ),
    .X(_2213_));
 sg13g2_nor2b_1 _3826_ (.A(net953),
    .B_N(net1053),
    .Y(_2214_));
 sg13g2_o21ai_1 _3827_ (.B1(net962),
    .Y(_2215_),
    .A1(_2213_),
    .A2(_2214_));
 sg13g2_nand3_1 _3828_ (.B(_2212_),
    .C(_2215_),
    .A(net1299),
    .Y(_2216_));
 sg13g2_o21ai_1 _3829_ (.B1(_2216_),
    .Y(_2217_),
    .A1(net1299),
    .A2(net349));
 sg13g2_inv_1 _3830_ (.Y(_0243_),
    .A(_2217_));
 sg13g2_nand2b_1 _3831_ (.Y(_2218_),
    .B(\s0.data_out[1][6] ),
    .A_N(net966));
 sg13g2_a21oi_1 _3832_ (.A1(_2140_),
    .A2(_2218_),
    .Y(_2219_),
    .B1(net964));
 sg13g2_nor2b_1 _3833_ (.A(net953),
    .B_N(net1049),
    .Y(_2220_));
 sg13g2_a21oi_1 _3834_ (.A1(net953),
    .A2(\s0.data_out[1][6] ),
    .Y(_2221_),
    .B1(_2220_));
 sg13g2_o21ai_1 _3835_ (.B1(net1299),
    .Y(_2222_),
    .A1(_2458_),
    .A2(_2221_));
 sg13g2_or2_1 _3836_ (.X(_2223_),
    .B(net491),
    .A(net1299));
 sg13g2_o21ai_1 _3837_ (.B1(_2223_),
    .Y(_2224_),
    .A1(_2219_),
    .A2(_2222_));
 sg13g2_inv_1 _3838_ (.Y(_0244_),
    .A(net492));
 sg13g2_nand2b_1 _3839_ (.Y(_2225_),
    .B(net495),
    .A_N(net966));
 sg13g2_a21oi_1 _3840_ (.A1(_2136_),
    .A2(_2225_),
    .Y(_2226_),
    .B1(net962));
 sg13g2_nor2b_1 _3841_ (.A(net953),
    .B_N(net1045),
    .Y(_2227_));
 sg13g2_a21oi_1 _3842_ (.A1(net954),
    .A2(net495),
    .Y(_2228_),
    .B1(_2227_));
 sg13g2_o21ai_1 _3843_ (.B1(net1298),
    .Y(_2229_),
    .A1(_2458_),
    .A2(_2228_));
 sg13g2_or2_1 _3844_ (.X(_2230_),
    .B(net553),
    .A(net1298));
 sg13g2_o21ai_1 _3845_ (.B1(_2230_),
    .Y(_2231_),
    .A1(_2226_),
    .A2(_2229_));
 sg13g2_inv_1 _3846_ (.Y(_0245_),
    .A(_2231_));
 sg13g2_mux2_1 _3847_ (.A0(\s0.data_out[2][2] ),
    .A1(\s0.data_out[1][2] ),
    .S(net955),
    .X(_2232_));
 sg13g2_a21o_1 _3848_ (.A2(_2232_),
    .A1(net949),
    .B1(_2192_),
    .X(_2233_));
 sg13g2_a21oi_1 _3849_ (.A1(net961),
    .A2(_2233_),
    .Y(_2234_),
    .B1(_2191_));
 sg13g2_or2_1 _3850_ (.X(_2235_),
    .B(_2234_),
    .A(net1268));
 sg13g2_mux2_1 _3851_ (.A0(\s0.data_out[2][1] ),
    .A1(\s0.data_out[1][1] ),
    .S(net955),
    .X(_2236_));
 sg13g2_a21oi_1 _3852_ (.A1(net949),
    .A2(_2236_),
    .Y(_2237_),
    .B1(_2186_));
 sg13g2_nand2b_1 _3853_ (.Y(_2238_),
    .B(net961),
    .A_N(_2237_));
 sg13g2_and2_1 _3854_ (.A(_2184_),
    .B(_2238_),
    .X(_2239_));
 sg13g2_mux2_1 _3855_ (.A0(\s0.data_out[2][0] ),
    .A1(\s0.data_out[1][0] ),
    .S(net955),
    .X(_2240_));
 sg13g2_a21oi_1 _3856_ (.A1(net950),
    .A2(_2240_),
    .Y(_2241_),
    .B1(_2179_));
 sg13g2_nand2b_1 _3857_ (.Y(_2242_),
    .B(net961),
    .A_N(_2241_));
 sg13g2_a221oi_1 _3858_ (.B2(_2177_),
    .C1(net1281),
    .B1(_2242_),
    .A1(net1273),
    .Y(_2243_),
    .A2(_2239_));
 sg13g2_o21ai_1 _3859_ (.B1(_2235_),
    .Y(_2244_),
    .A1(net1273),
    .A2(_2239_));
 sg13g2_nand2_1 _3860_ (.Y(_2245_),
    .A(net955),
    .B(net513));
 sg13g2_mux2_1 _3861_ (.A0(\s0.data_out[2][3] ),
    .A1(\s0.data_out[1][3] ),
    .S(net958),
    .X(_2246_));
 sg13g2_a21oi_1 _3862_ (.A1(net950),
    .A2(_2246_),
    .Y(_2247_),
    .B1(_2200_));
 sg13g2_nand2b_1 _3863_ (.Y(_2248_),
    .B(net961),
    .A_N(_2247_));
 sg13g2_and2_1 _3864_ (.A(_2198_),
    .B(_2248_),
    .X(_2249_));
 sg13g2_a22oi_1 _3865_ (.Y(_2250_),
    .B1(_2249_),
    .B2(net1261),
    .A2(_2234_),
    .A1(net1268));
 sg13g2_o21ai_1 _3866_ (.B1(_2250_),
    .Y(_2251_),
    .A1(_2243_),
    .A2(_2244_));
 sg13g2_nand2_1 _3867_ (.Y(_2252_),
    .A(net956),
    .B(net495));
 sg13g2_mux2_1 _3868_ (.A0(\s0.data_out[2][7] ),
    .A1(\s0.data_out[1][7] ),
    .S(net957),
    .X(_2253_));
 sg13g2_a21o_1 _3869_ (.A2(_2253_),
    .A1(net954),
    .B1(_2227_),
    .X(_2254_));
 sg13g2_a21oi_1 _3870_ (.A1(net964),
    .A2(_2254_),
    .Y(_2255_),
    .B1(_2226_));
 sg13g2_nand2_1 _3871_ (.Y(_2256_),
    .A(net956),
    .B(net590));
 sg13g2_mux2_1 _3872_ (.A0(\s0.data_out[2][6] ),
    .A1(\s0.data_out[1][6] ),
    .S(net957),
    .X(_2257_));
 sg13g2_a21o_1 _3873_ (.A2(_2257_),
    .A1(net954),
    .B1(_2220_),
    .X(_2258_));
 sg13g2_a21oi_1 _3874_ (.A1(net962),
    .A2(_2258_),
    .Y(_2259_),
    .B1(_2219_));
 sg13g2_a22oi_1 _3875_ (.Y(_2260_),
    .B1(_2259_),
    .B2(net1239),
    .A2(_2255_),
    .A1(net1232));
 sg13g2_or2_1 _3876_ (.X(_2261_),
    .B(_2255_),
    .A(net1232));
 sg13g2_or2_1 _3877_ (.X(_2262_),
    .B(_2259_),
    .A(net1239));
 sg13g2_nand3_1 _3878_ (.B(_2261_),
    .C(_2262_),
    .A(_2260_),
    .Y(_2263_));
 sg13g2_inv_1 _3879_ (.Y(_2264_),
    .A(_2263_));
 sg13g2_mux2_1 _3880_ (.A0(\s0.data_out[2][4] ),
    .A1(\s0.data_out[1][4] ),
    .S(net958),
    .X(_2265_));
 sg13g2_a21oi_1 _3881_ (.A1(net950),
    .A2(_2265_),
    .Y(_2266_),
    .B1(_2207_));
 sg13g2_o21ai_1 _3882_ (.B1(_2205_),
    .Y(_2267_),
    .A1(net930),
    .A2(_2266_));
 sg13g2_or2_1 _3883_ (.X(_2268_),
    .B(_2267_),
    .A(net1214));
 sg13g2_mux2_1 _3884_ (.A0(\s0.data_out[2][5] ),
    .A1(\s0.data_out[1][5] ),
    .S(net957),
    .X(_2269_));
 sg13g2_a21oi_1 _3885_ (.A1(net953),
    .A2(_2269_),
    .Y(_2270_),
    .B1(_2214_));
 sg13g2_nand2b_1 _3886_ (.Y(_2271_),
    .B(net962),
    .A_N(_2270_));
 sg13g2_nand3_1 _3887_ (.B(_2212_),
    .C(_2271_),
    .A(net1247),
    .Y(_2272_));
 sg13g2_nor2_1 _3888_ (.A(net1261),
    .B(_2249_),
    .Y(_2273_));
 sg13g2_a21oi_1 _3889_ (.A1(_2212_),
    .A2(_2271_),
    .Y(_2274_),
    .B1(net1247));
 sg13g2_xnor2_1 _3890_ (.Y(_2275_),
    .A(net1214),
    .B(_2267_));
 sg13g2_nor3_1 _3891_ (.A(_2273_),
    .B(_2274_),
    .C(_2275_),
    .Y(_2276_));
 sg13g2_nand4_1 _3892_ (.B(_2264_),
    .C(_2272_),
    .A(_2251_),
    .Y(_2277_),
    .D(_2276_));
 sg13g2_o21ai_1 _3893_ (.B1(_2272_),
    .Y(_2278_),
    .A1(_2268_),
    .A2(_2274_));
 sg13g2_nor2b_1 _3894_ (.A(_2263_),
    .B_N(_2278_),
    .Y(_2279_));
 sg13g2_nor2b_1 _3895_ (.A(_2260_),
    .B_N(_2261_),
    .Y(_2280_));
 sg13g2_nor3_1 _3896_ (.A(_2170_),
    .B(_2279_),
    .C(_2280_),
    .Y(_2281_));
 sg13g2_or2_1 _3897_ (.X(_2282_),
    .B(net1208),
    .A(net300));
 sg13g2_a21oi_1 _3898_ (.A1(_2277_),
    .A2(_2281_),
    .Y(_0246_),
    .B1(_2282_));
 sg13g2_and2_1 _3899_ (.A(net1291),
    .B(net306),
    .X(_0247_));
 sg13g2_o21ai_1 _3900_ (.B1(net952),
    .Y(_2283_),
    .A1(net1225),
    .A2(net943));
 sg13g2_a21oi_1 _3901_ (.A1(net1222),
    .A2(net947),
    .Y(_2284_),
    .B1(_2283_));
 sg13g2_a21oi_1 _3902_ (.A1(net928),
    .A2(_2167_),
    .Y(_2285_),
    .B1(_2284_));
 sg13g2_o21ai_1 _3903_ (.B1(_2284_),
    .Y(_2286_),
    .A1(\s0.was_valid_out[0] [0]),
    .A2(net947));
 sg13g2_nor2_1 _3904_ (.A(net943),
    .B(_2283_),
    .Y(_2287_));
 sg13g2_o21ai_1 _3905_ (.B1(net929),
    .Y(_2288_),
    .A1(\s0.was_valid_out[0] [0]),
    .A2(net956));
 sg13g2_nand2_1 _3906_ (.Y(_2289_),
    .A(_2286_),
    .B(_2288_));
 sg13g2_o21ai_1 _3907_ (.B1(net1298),
    .Y(_2290_),
    .A1(_2287_),
    .A2(_2289_));
 sg13g2_a21oi_1 _3908_ (.A1(_2442_),
    .A2(_2285_),
    .Y(_0248_),
    .B1(_2290_));
 sg13g2_and2_1 _3909_ (.A(net1299),
    .B(_2285_),
    .X(_0249_));
 sg13g2_mux2_1 _3910_ (.A0(\s0.data_out[0][0] ),
    .A1(\s0.data_out[1][0] ),
    .S(net955),
    .X(_2291_));
 sg13g2_nand2_1 _3911_ (.Y(_2292_),
    .A(net928),
    .B(_2291_));
 sg13g2_and2_1 _3912_ (.A(net941),
    .B(\s0.data_out[0][0] ),
    .X(_2293_));
 sg13g2_nor2b_1 _3913_ (.A(net940),
    .B_N(net1073),
    .Y(_2294_));
 sg13g2_o21ai_1 _3914_ (.B1(net951),
    .Y(_2295_),
    .A1(_2293_),
    .A2(_2294_));
 sg13g2_nand3_1 _3915_ (.B(_2292_),
    .C(_2295_),
    .A(net1293),
    .Y(_2296_));
 sg13g2_o21ai_1 _3916_ (.B1(_2296_),
    .Y(_2297_),
    .A1(net1293),
    .A2(net448));
 sg13g2_inv_1 _3917_ (.Y(_0250_),
    .A(net449));
 sg13g2_mux2_1 _3918_ (.A0(\s0.data_out[0][1] ),
    .A1(\s0.data_out[1][1] ),
    .S(net955),
    .X(_2298_));
 sg13g2_nand2_1 _3919_ (.Y(_2299_),
    .A(net928),
    .B(_2298_));
 sg13g2_and2_1 _3920_ (.A(net942),
    .B(\s0.data_out[0][1] ),
    .X(_2300_));
 sg13g2_nor2b_1 _3921_ (.A(net942),
    .B_N(net1069),
    .Y(_2301_));
 sg13g2_o21ai_1 _3922_ (.B1(net951),
    .Y(_2302_),
    .A1(_2300_),
    .A2(_2301_));
 sg13g2_nand3_1 _3923_ (.B(_2299_),
    .C(_2302_),
    .A(net1293),
    .Y(_2303_));
 sg13g2_o21ai_1 _3924_ (.B1(_2303_),
    .Y(_2304_),
    .A1(net1293),
    .A2(net396));
 sg13g2_inv_1 _3925_ (.Y(_0251_),
    .A(net397));
 sg13g2_mux2_1 _3926_ (.A0(\s0.data_out[0][2] ),
    .A1(\s0.data_out[1][2] ),
    .S(net955),
    .X(_2305_));
 sg13g2_nand2_1 _3927_ (.Y(_2306_),
    .A(net928),
    .B(_2305_));
 sg13g2_and2_1 _3928_ (.A(net940),
    .B(\s0.data_out[0][2] ),
    .X(_2307_));
 sg13g2_nor2b_1 _3929_ (.A(net942),
    .B_N(net1065),
    .Y(_2308_));
 sg13g2_o21ai_1 _3930_ (.B1(net951),
    .Y(_2309_),
    .A1(_2307_),
    .A2(_2308_));
 sg13g2_nand3_1 _3931_ (.B(_2306_),
    .C(_2309_),
    .A(net1292),
    .Y(_2310_));
 sg13g2_o21ai_1 _3932_ (.B1(_2310_),
    .Y(_2311_),
    .A1(net1293),
    .A2(net458));
 sg13g2_inv_1 _3933_ (.Y(_0252_),
    .A(net459));
 sg13g2_nand2b_1 _3934_ (.Y(_2312_),
    .B(net348),
    .A_N(net955));
 sg13g2_a21oi_1 _3935_ (.A1(_2245_),
    .A2(_2312_),
    .Y(_2313_),
    .B1(net951));
 sg13g2_nor2b_1 _3936_ (.A(net941),
    .B_N(net1061),
    .Y(_2314_));
 sg13g2_a21oi_1 _3937_ (.A1(net941),
    .A2(net348),
    .Y(_2315_),
    .B1(_2314_));
 sg13g2_o21ai_1 _3938_ (.B1(net1293),
    .Y(_2316_),
    .A1(net928),
    .A2(_2315_));
 sg13g2_or2_1 _3939_ (.X(_2317_),
    .B(net513),
    .A(net1293));
 sg13g2_o21ai_1 _3940_ (.B1(_2317_),
    .Y(_2318_),
    .A1(_2313_),
    .A2(_2316_));
 sg13g2_inv_1 _3941_ (.Y(_0253_),
    .A(net514));
 sg13g2_mux2_1 _3942_ (.A0(\s0.data_out[0][4] ),
    .A1(\s0.data_out[1][4] ),
    .S(net956),
    .X(_2319_));
 sg13g2_nand2_1 _3943_ (.Y(_2320_),
    .A(net929),
    .B(_2319_));
 sg13g2_and2_1 _3944_ (.A(net945),
    .B(\s0.data_out[0][4] ),
    .X(_2321_));
 sg13g2_nor2b_1 _3945_ (.A(net942),
    .B_N(net1057),
    .Y(_2322_));
 sg13g2_o21ai_1 _3946_ (.B1(net952),
    .Y(_2323_),
    .A1(_2321_),
    .A2(_2322_));
 sg13g2_nand3_1 _3947_ (.B(_2320_),
    .C(_2323_),
    .A(net1298),
    .Y(_2324_));
 sg13g2_o21ai_1 _3948_ (.B1(_2324_),
    .Y(_2325_),
    .A1(net1298),
    .A2(net394));
 sg13g2_inv_1 _3949_ (.Y(_0254_),
    .A(_2325_));
 sg13g2_mux2_1 _3950_ (.A0(\s0.data_out[0][5] ),
    .A1(\s0.data_out[1][5] ),
    .S(net956),
    .X(_2326_));
 sg13g2_nand2_1 _3951_ (.Y(_2327_),
    .A(net929),
    .B(_2326_));
 sg13g2_and2_1 _3952_ (.A(net944),
    .B(\s0.data_out[0][5] ),
    .X(_2328_));
 sg13g2_nor2b_1 _3953_ (.A(net943),
    .B_N(net1053),
    .Y(_2329_));
 sg13g2_o21ai_1 _3954_ (.B1(net952),
    .Y(_2330_),
    .A1(_2328_),
    .A2(_2329_));
 sg13g2_nand3_1 _3955_ (.B(_2327_),
    .C(_2330_),
    .A(net1295),
    .Y(_2331_));
 sg13g2_o21ai_1 _3956_ (.B1(_2331_),
    .Y(_2332_),
    .A1(net1295),
    .A2(net479));
 sg13g2_inv_1 _3957_ (.Y(_0255_),
    .A(_2332_));
 sg13g2_nand2b_1 _3958_ (.Y(_2333_),
    .B(net351),
    .A_N(net956));
 sg13g2_a21oi_1 _3959_ (.A1(_2256_),
    .A2(_2333_),
    .Y(_2334_),
    .B1(net952));
 sg13g2_nor2b_1 _3960_ (.A(net945),
    .B_N(net1049),
    .Y(_2335_));
 sg13g2_a21oi_1 _3961_ (.A1(net943),
    .A2(net351),
    .Y(_2336_),
    .B1(_2335_));
 sg13g2_o21ai_1 _3962_ (.B1(net1295),
    .Y(_2337_),
    .A1(net929),
    .A2(_2336_));
 sg13g2_or2_1 _3963_ (.X(_2338_),
    .B(net590),
    .A(net1295));
 sg13g2_o21ai_1 _3964_ (.B1(_2338_),
    .Y(_2339_),
    .A1(_2334_),
    .A2(_2337_));
 sg13g2_inv_1 _3965_ (.Y(_0256_),
    .A(_2339_));
 sg13g2_nand2b_1 _3966_ (.Y(_2340_),
    .B(net334),
    .A_N(net956));
 sg13g2_a21oi_1 _3967_ (.A1(_2252_),
    .A2(_2340_),
    .Y(_2341_),
    .B1(net952));
 sg13g2_nor2b_1 _3968_ (.A(net944),
    .B_N(net1045),
    .Y(_2342_));
 sg13g2_a21oi_1 _3969_ (.A1(net945),
    .A2(net334),
    .Y(_2343_),
    .B1(_2342_));
 sg13g2_o21ai_1 _3970_ (.B1(net1295),
    .Y(_2344_),
    .A1(net929),
    .A2(_2343_));
 sg13g2_or2_1 _3971_ (.X(_2345_),
    .B(net495),
    .A(net1299));
 sg13g2_o21ai_1 _3972_ (.B1(_2345_),
    .Y(_2346_),
    .A1(_2341_),
    .A2(_2344_));
 sg13g2_inv_1 _3973_ (.Y(_0257_),
    .A(_2346_));
 sg13g2_nand2_1 _3974_ (.Y(_2347_),
    .A(net946),
    .B(net345));
 sg13g2_o21ai_1 _3975_ (.B1(_2347_),
    .Y(_2348_),
    .A1(net946),
    .A2(_2493_));
 sg13g2_a21oi_1 _3976_ (.A1(net942),
    .A2(_2348_),
    .Y(_2349_),
    .B1(_2308_));
 sg13g2_o21ai_1 _3977_ (.B1(_2306_),
    .Y(_2350_),
    .A1(net928),
    .A2(_2349_));
 sg13g2_mux2_1 _3978_ (.A0(\s0.data_out[1][1] ),
    .A1(\s0.data_out[0][1] ),
    .S(net948),
    .X(_2351_));
 sg13g2_a21oi_1 _3979_ (.A1(net942),
    .A2(_2351_),
    .Y(_2352_),
    .B1(_2301_));
 sg13g2_nand2b_1 _3980_ (.Y(_2353_),
    .B(net951),
    .A_N(_2352_));
 sg13g2_nand3_1 _3981_ (.B(_2299_),
    .C(_2353_),
    .A(net1274),
    .Y(_2354_));
 sg13g2_mux2_1 _3982_ (.A0(\s0.data_out[1][0] ),
    .A1(\s0.data_out[0][0] ),
    .S(net946),
    .X(_2355_));
 sg13g2_a21oi_1 _3983_ (.A1(net942),
    .A2(_2355_),
    .Y(_2356_),
    .B1(_2294_));
 sg13g2_o21ai_1 _3984_ (.B1(_2292_),
    .Y(_2357_),
    .A1(net928),
    .A2(_2356_));
 sg13g2_nor2b_1 _3985_ (.A(net1281),
    .B_N(_2357_),
    .Y(_2358_));
 sg13g2_a21oi_1 _3986_ (.A1(_2299_),
    .A2(_2353_),
    .Y(_2359_),
    .B1(net1274));
 sg13g2_a221oi_1 _3987_ (.B2(_2358_),
    .C1(_2359_),
    .B1(_2354_),
    .A1(net1211),
    .Y(_2360_),
    .A2(_2350_));
 sg13g2_nand2_1 _3988_ (.Y(_2361_),
    .A(net946),
    .B(net348));
 sg13g2_nand2b_1 _3989_ (.Y(_2362_),
    .B(\s0.data_out[1][3] ),
    .A_N(net946));
 sg13g2_a21oi_1 _3990_ (.A1(_2361_),
    .A2(_2362_),
    .Y(_2363_),
    .B1(_2465_));
 sg13g2_or2_1 _3991_ (.X(_2364_),
    .B(_2363_),
    .A(_2314_));
 sg13g2_a21oi_1 _3992_ (.A1(net951),
    .A2(_2364_),
    .Y(_2365_),
    .B1(_2313_));
 sg13g2_and2_1 _3993_ (.A(net1261),
    .B(_2365_),
    .X(_2366_));
 sg13g2_nor2_1 _3994_ (.A(net1211),
    .B(_2350_),
    .Y(_2367_));
 sg13g2_or3_1 _3995_ (.A(_2360_),
    .B(_2366_),
    .C(_2367_),
    .X(_2368_));
 sg13g2_mux2_1 _3996_ (.A0(\s0.data_out[1][7] ),
    .A1(\s0.data_out[0][7] ),
    .S(net948),
    .X(_2369_));
 sg13g2_a21o_1 _3997_ (.A2(_2369_),
    .A1(net943),
    .B1(_2342_),
    .X(_2370_));
 sg13g2_a21oi_1 _3998_ (.A1(net954),
    .A2(_2370_),
    .Y(_2371_),
    .B1(_2341_));
 sg13g2_mux2_1 _3999_ (.A0(\s0.data_out[1][6] ),
    .A1(\s0.data_out[0][6] ),
    .S(net947),
    .X(_2372_));
 sg13g2_a21o_1 _4000_ (.A2(_2372_),
    .A1(net943),
    .B1(_2335_),
    .X(_2373_));
 sg13g2_a21oi_1 _4001_ (.A1(net952),
    .A2(_2373_),
    .Y(_2374_),
    .B1(_2334_));
 sg13g2_a22oi_1 _4002_ (.Y(_2375_),
    .B1(_2374_),
    .B2(net1241),
    .A2(_2371_),
    .A1(net1232));
 sg13g2_or2_1 _4003_ (.X(_2376_),
    .B(_2374_),
    .A(net1241));
 sg13g2_or2_1 _4004_ (.X(_2377_),
    .B(_2371_),
    .A(net1232));
 sg13g2_inv_1 _4005_ (.Y(_2378_),
    .A(_2377_));
 sg13g2_and3_1 _4006_ (.X(_2379_),
    .A(_2375_),
    .B(_2376_),
    .C(_2377_));
 sg13g2_mux2_1 _4007_ (.A0(\s0.data_out[1][4] ),
    .A1(\s0.data_out[0][4] ),
    .S(net948),
    .X(_2380_));
 sg13g2_a21oi_1 _4008_ (.A1(net943),
    .A2(_2380_),
    .Y(_2381_),
    .B1(_2322_));
 sg13g2_o21ai_1 _4009_ (.B1(_2320_),
    .Y(_2382_),
    .A1(net928),
    .A2(_2381_));
 sg13g2_or2_1 _4010_ (.X(_2383_),
    .B(_2382_),
    .A(net1214));
 sg13g2_mux2_1 _4011_ (.A0(\s0.data_out[1][5] ),
    .A1(\s0.data_out[0][5] ),
    .S(net947),
    .X(_2384_));
 sg13g2_a21oi_1 _4012_ (.A1(net943),
    .A2(_2384_),
    .Y(_2385_),
    .B1(_2329_));
 sg13g2_nand2b_1 _4013_ (.Y(_2386_),
    .B(net952),
    .A_N(_2385_));
 sg13g2_and2_1 _4014_ (.A(_2327_),
    .B(_2386_),
    .X(_2387_));
 sg13g2_nand2_1 _4015_ (.Y(_2388_),
    .A(net1247),
    .B(_2387_));
 sg13g2_or2_1 _4016_ (.X(_2389_),
    .B(_2365_),
    .A(net1261));
 sg13g2_nor2_1 _4017_ (.A(net1247),
    .B(_2387_),
    .Y(_2390_));
 sg13g2_xnor2_1 _4018_ (.Y(_2391_),
    .A(net1254),
    .B(_2382_));
 sg13g2_xor2_1 _4019_ (.B(_2387_),
    .A(net1247),
    .X(_2392_));
 sg13g2_and4_1 _4020_ (.A(_2379_),
    .B(_2389_),
    .C(_2391_),
    .D(_2392_),
    .X(_2393_));
 sg13g2_o21ai_1 _4021_ (.B1(_2388_),
    .Y(_2394_),
    .A1(_2383_),
    .A2(_2390_));
 sg13g2_o21ai_1 _4022_ (.B1(_2285_),
    .Y(_2395_),
    .A1(_2375_),
    .A2(_2378_));
 sg13g2_a221oi_1 _4023_ (.B2(_2379_),
    .C1(_2395_),
    .B1(_2394_),
    .A1(_2368_),
    .Y(_2396_),
    .A2(_2393_));
 sg13g2_nor3_1 _4024_ (.A(net297),
    .B(net1208),
    .C(_2396_),
    .Y(_0258_));
 sg13g2_and2_1 _4025_ (.A(net1289),
    .B(net305),
    .X(_0259_));
 sg13g2_a21oi_1 _4026_ (.A1(net363),
    .A2(_2465_),
    .Y(_2397_),
    .B1(net1225));
 sg13g2_o21ai_1 _4027_ (.B1(net1294),
    .Y(_2398_),
    .A1(net947),
    .A2(net944));
 sg13g2_nor2_1 _4028_ (.A(_2397_),
    .B(_2398_),
    .Y(_0260_));
 sg13g2_nor2_1 _4029_ (.A(net1225),
    .B(_2398_),
    .Y(_0261_));
 sg13g2_a21oi_1 _4030_ (.A1(net946),
    .A2(net377),
    .Y(_2399_),
    .B1(net940));
 sg13g2_nor2b_1 _4031_ (.A(net1073),
    .B_N(net940),
    .Y(_2400_));
 sg13g2_nor3_1 _4032_ (.A(net1218),
    .B(_2399_),
    .C(_2400_),
    .Y(_2401_));
 sg13g2_a21o_1 _4033_ (.A2(net377),
    .A1(net1218),
    .B1(_2401_),
    .X(_0262_));
 sg13g2_a21oi_1 _4034_ (.A1(net946),
    .A2(net392),
    .Y(_2402_),
    .B1(net940));
 sg13g2_nor2b_1 _4035_ (.A(net1069),
    .B_N(net940),
    .Y(_2403_));
 sg13g2_o21ai_1 _4036_ (.B1(net1292),
    .Y(_2404_),
    .A1(_2402_),
    .A2(_2403_));
 sg13g2_o21ai_1 _4037_ (.B1(_2404_),
    .Y(_2405_),
    .A1(net1292),
    .A2(net392));
 sg13g2_inv_1 _4038_ (.Y(_0263_),
    .A(_2405_));
 sg13g2_nor2_1 _4039_ (.A(net1292),
    .B(net345),
    .Y(_2406_));
 sg13g2_nand2_1 _4040_ (.Y(_2407_),
    .A(net940),
    .B(net1065));
 sg13g2_o21ai_1 _4041_ (.B1(_2407_),
    .Y(_2408_),
    .A1(net940),
    .A2(_2347_));
 sg13g2_inv_1 _4042_ (.Y(_2409_),
    .A(_2408_));
 sg13g2_a21oi_1 _4043_ (.A1(net1292),
    .A2(_2409_),
    .Y(_0264_),
    .B1(_2406_));
 sg13g2_nor2_1 _4044_ (.A(net1292),
    .B(net348),
    .Y(_2410_));
 sg13g2_nor2_1 _4045_ (.A(net941),
    .B(_2361_),
    .Y(_2411_));
 sg13g2_a21oi_1 _4046_ (.A1(net941),
    .A2(net1061),
    .Y(_2412_),
    .B1(_2411_));
 sg13g2_a21oi_1 _4047_ (.A1(net1292),
    .A2(_2412_),
    .Y(_0265_),
    .B1(_2410_));
 sg13g2_a21o_1 _4048_ (.A2(net374),
    .A1(net946),
    .B1(net941),
    .X(_2413_));
 sg13g2_o21ai_1 _4049_ (.B1(_2413_),
    .Y(_2414_),
    .A1(_2465_),
    .A2(net1057));
 sg13g2_nor2_1 _4050_ (.A(net1218),
    .B(_2414_),
    .Y(_2415_));
 sg13g2_a21oi_1 _4051_ (.A1(net1218),
    .A2(net374),
    .Y(_2416_),
    .B1(_2415_));
 sg13g2_inv_1 _4052_ (.Y(_0266_),
    .A(_2416_));
 sg13g2_nor2_1 _4053_ (.A(net1294),
    .B(net344),
    .Y(_2417_));
 sg13g2_a21o_1 _4054_ (.A2(net344),
    .A1(net947),
    .B1(net944),
    .X(_2418_));
 sg13g2_o21ai_1 _4055_ (.B1(_2418_),
    .Y(_2419_),
    .A1(_2465_),
    .A2(net1053));
 sg13g2_a21oi_1 _4056_ (.A1(net1294),
    .A2(_2419_),
    .Y(_0267_),
    .B1(_2417_));
 sg13g2_nor2_1 _4057_ (.A(net1294),
    .B(net351),
    .Y(_2420_));
 sg13g2_a21o_1 _4058_ (.A2(net351),
    .A1(net947),
    .B1(net944),
    .X(_2421_));
 sg13g2_o21ai_1 _4059_ (.B1(_2421_),
    .Y(_2422_),
    .A1(_2465_),
    .A2(net1049));
 sg13g2_a21oi_1 _4060_ (.A1(net1294),
    .A2(_2422_),
    .Y(_0268_),
    .B1(_2420_));
 sg13g2_nor2_1 _4061_ (.A(net1294),
    .B(net334),
    .Y(_2423_));
 sg13g2_a21o_1 _4062_ (.A2(net334),
    .A1(net947),
    .B1(net944),
    .X(_2424_));
 sg13g2_o21ai_1 _4063_ (.B1(_2424_),
    .Y(_2425_),
    .A1(_2465_),
    .A2(net1045));
 sg13g2_a21oi_1 _4064_ (.A1(net1294),
    .A2(_2425_),
    .Y(_0269_),
    .B1(_2423_));
 sg13g2_or2_1 _4065_ (.X(_2426_),
    .B(_2419_),
    .A(net1246));
 sg13g2_a22oi_1 _4066_ (.Y(_2427_),
    .B1(_2419_),
    .B2(net1246),
    .A2(_2414_),
    .A1(net1254));
 sg13g2_o21ai_1 _4067_ (.B1(net1274),
    .Y(_2428_),
    .A1(_2402_),
    .A2(_2403_));
 sg13g2_nor3_1 _4068_ (.A(net1281),
    .B(_2399_),
    .C(_2400_),
    .Y(_2429_));
 sg13g2_nor3_1 _4069_ (.A(net1274),
    .B(_2402_),
    .C(_2403_),
    .Y(_2430_));
 sg13g2_a221oi_1 _4070_ (.B2(_2429_),
    .C1(_2430_),
    .B1(_2428_),
    .A1(net1211),
    .Y(_2431_),
    .A2(_2408_));
 sg13g2_a221oi_1 _4071_ (.B2(net1260),
    .C1(_2431_),
    .B1(_2412_),
    .A1(net1268),
    .Y(_2432_),
    .A2(_2409_));
 sg13g2_nand2b_1 _4072_ (.Y(_2433_),
    .B(net1214),
    .A_N(_2414_));
 sg13g2_o21ai_1 _4073_ (.B1(_2433_),
    .Y(_2434_),
    .A1(net1260),
    .A2(_2412_));
 sg13g2_o21ai_1 _4074_ (.B1(_2427_),
    .Y(_2435_),
    .A1(_2432_),
    .A2(_2434_));
 sg13g2_a22oi_1 _4075_ (.Y(_2436_),
    .B1(_2426_),
    .B2(_2435_),
    .A2(_2422_),
    .A1(net1241));
 sg13g2_nand2b_1 _4076_ (.Y(_2437_),
    .B(_2474_),
    .A_N(_2422_));
 sg13g2_o21ai_1 _4077_ (.B1(_2437_),
    .Y(_2438_),
    .A1(net1232),
    .A2(_2425_));
 sg13g2_a21oi_1 _4078_ (.A1(net1232),
    .A2(_2425_),
    .Y(_2439_),
    .B1(net1227));
 sg13g2_o21ai_1 _4079_ (.B1(_2439_),
    .Y(_2440_),
    .A1(_2436_),
    .A2(_2438_));
 sg13g2_nor2_1 _4080_ (.A(net312),
    .B(net1208),
    .Y(_2441_));
 sg13g2_and2_1 _4081_ (.A(_2440_),
    .B(_2441_),
    .X(_0270_));
 sg13g2_and2_1 _4082_ (.A(net1342),
    .B(net314),
    .X(_0271_));
 sg13g2_inv_1 _4083_ (.Y(_2442_),
    .A(net328));
 sg13g2_inv_1 _4084_ (.Y(_2443_),
    .A(net319));
 sg13g2_inv_1 _4085_ (.Y(_2444_),
    .A(net326));
 sg13g2_inv_1 _4086_ (.Y(_2445_),
    .A(net346));
 sg13g2_inv_1 _4087_ (.Y(_2446_),
    .A(net321));
 sg13g2_inv_1 _4088_ (.Y(_2447_),
    .A(net323));
 sg13g2_inv_1 _4089_ (.Y(_2448_),
    .A(net1093));
 sg13g2_inv_4 _4090_ (.A(net1228),
    .Y(_2449_));
 sg13g2_inv_4 _4091_ (.A(net1337),
    .Y(_2450_));
 sg13g2_inv_1 _4092_ (.Y(_2451_),
    .A(net1105));
 sg13g2_inv_1 _4093_ (.Y(_2452_),
    .A(net1128));
 sg13g2_inv_1 _4094_ (.Y(_2453_),
    .A(net1118));
 sg13g2_inv_1 _4095_ (.Y(_2454_),
    .A(net1082));
 sg13g2_inv_1 _4096_ (.Y(_2455_),
    .A(net973));
 sg13g2_inv_2 _4097_ (.Y(_2456_),
    .A(net1194));
 sg13g2_inv_1 _4098_ (.Y(_2457_),
    .A(net1203));
 sg13g2_inv_2 _4099_ (.Y(_2458_),
    .A(net962));
 sg13g2_inv_1 _4100_ (.Y(_2459_),
    .A(net952));
 sg13g2_inv_1 _4101_ (.Y(_2460_),
    .A(net1181));
 sg13g2_inv_2 _4102_ (.Y(_2461_),
    .A(net1171));
 sg13g2_inv_2 _4103_ (.Y(_2462_),
    .A(net1160));
 sg13g2_inv_1 _4104_ (.Y(_2463_),
    .A(net1148));
 sg13g2_inv_2 _4105_ (.Y(_2464_),
    .A(net1138));
 sg13g2_inv_2 _4106_ (.Y(_2465_),
    .A(net944));
 sg13g2_inv_1 _4107_ (.Y(_2466_),
    .A(net1037));
 sg13g2_inv_1 _4108_ (.Y(_2467_),
    .A(net1025));
 sg13g2_inv_2 _4109_ (.Y(_2468_),
    .A(net1012));
 sg13g2_inv_1 _4110_ (.Y(_2469_),
    .A(net1004));
 sg13g2_inv_1 _4111_ (.Y(_2470_),
    .A(net994));
 sg13g2_inv_2 _4112_ (.Y(_2471_),
    .A(net983));
 sg13g2_inv_1 _4113_ (.Y(_2472_),
    .A(net364));
 sg13g2_inv_1 _4114_ (.Y(_2473_),
    .A(net356));
 sg13g2_inv_2 _4115_ (.Y(_2474_),
    .A(net1239));
 sg13g2_inv_1 _4116_ (.Y(_2475_),
    .A(net361));
 sg13g2_inv_1 _4117_ (.Y(_2476_),
    .A(net1254));
 sg13g2_inv_1 _4118_ (.Y(_2477_),
    .A(net359));
 sg13g2_inv_1 _4119_ (.Y(_2478_),
    .A(net366));
 sg13g2_inv_1 _4120_ (.Y(_2479_),
    .A(\s0.data_out[21][2] ));
 sg13g2_inv_2 _4121_ (.Y(_2480_),
    .A(net1268));
 sg13g2_inv_1 _4122_ (.Y(_2481_),
    .A(\s0.data_out[21][1] ));
 sg13g2_inv_1 _4123_ (.Y(_2482_),
    .A(net368));
 sg13g2_inv_1 _4124_ (.Y(_2483_),
    .A(\s0.data_out[19][2] ));
 sg13g2_inv_2 _4125_ (.Y(_2484_),
    .A(net493));
 sg13g2_inv_2 _4126_ (.Y(_2485_),
    .A(net550));
 sg13g2_inv_1 _4127_ (.Y(_2486_),
    .A(net386));
 sg13g2_inv_1 _4128_ (.Y(_2487_),
    .A(\s0.data_out[13][2] ));
 sg13g2_inv_1 _4129_ (.Y(_2488_),
    .A(\s0.data_out[12][3] ));
 sg13g2_inv_1 _4130_ (.Y(_2489_),
    .A(\s0.data_out[9][2] ));
 sg13g2_inv_2 _4131_ (.Y(_2490_),
    .A(\s0.data_out[9][5] ));
 sg13g2_inv_1 _4132_ (.Y(_2491_),
    .A(\s0.data_out[7][2] ));
 sg13g2_inv_1 _4133_ (.Y(_2492_),
    .A(\s0.data_out[3][2] ));
 sg13g2_inv_1 _4134_ (.Y(_2493_),
    .A(\s0.data_out[1][2] ));
 sg13g2_nor2_1 _4135_ (.A(\s0.was_valid_out[21] [0]),
    .B(net1204),
    .Y(_2494_));
 sg13g2_nand2_1 _4136_ (.Y(_2495_),
    .A(net1281),
    .B(net913));
 sg13g2_o21ai_1 _4137_ (.B1(_2495_),
    .Y(net2),
    .A1(_2482_),
    .A2(net913));
 sg13g2_nand2_1 _4138_ (.Y(_2496_),
    .A(net1273),
    .B(net913));
 sg13g2_o21ai_1 _4139_ (.B1(_2496_),
    .Y(net3),
    .A1(_2481_),
    .A2(net913));
 sg13g2_nor2_1 _4140_ (.A(\s0.data_out[21][2] ),
    .B(net913),
    .Y(_2497_));
 sg13g2_a21oi_1 _4141_ (.A1(net1211),
    .A2(net913),
    .Y(net4),
    .B1(_2497_));
 sg13g2_nand2_1 _4142_ (.Y(_2498_),
    .A(net1260),
    .B(net912));
 sg13g2_o21ai_1 _4143_ (.B1(_2498_),
    .Y(net5),
    .A1(_2478_),
    .A2(net913));
 sg13g2_nor2_1 _4144_ (.A(\s0.data_out[21][4] ),
    .B(net912),
    .Y(_2499_));
 sg13g2_a21oi_1 _4145_ (.A1(net1214),
    .A2(net912),
    .Y(net6),
    .B1(_2499_));
 sg13g2_nand2_1 _4146_ (.Y(_2500_),
    .A(net1246),
    .B(net912));
 sg13g2_o21ai_1 _4147_ (.B1(_2500_),
    .Y(net7),
    .A1(_2475_),
    .A2(net912));
 sg13g2_nor2_1 _4148_ (.A(\s0.data_out[21][6] ),
    .B(net912),
    .Y(_2501_));
 sg13g2_a21oi_1 _4149_ (.A1(_2474_),
    .A2(net912),
    .Y(net8),
    .B1(_2501_));
 sg13g2_nand2_1 _4150_ (.Y(_2502_),
    .A(net1231),
    .B(_2494_));
 sg13g2_o21ai_1 _4151_ (.B1(_2502_),
    .Y(net9),
    .A1(_2472_),
    .A2(net912));
 sg13g2_and2_1 _4152_ (.A(net1294),
    .B(net312),
    .X(_0000_));
 sg13g2_o21ai_1 _4153_ (.B1(net1204),
    .Y(_2503_),
    .A1(net1225),
    .A2(net1195));
 sg13g2_nor2b_1 _4154_ (.A(net1225),
    .B_N(net1200),
    .Y(_2504_));
 sg13g2_or2_1 _4155_ (.X(_2505_),
    .B(_2504_),
    .A(_2503_));
 sg13g2_nor2b_1 _4156_ (.A(net1225),
    .B_N(net1207),
    .Y(_2506_));
 sg13g2_o21ai_1 _4157_ (.B1(_2505_),
    .Y(_2507_),
    .A1(net1205),
    .A2(_2506_));
 sg13g2_nor2_1 _4158_ (.A(\s0.was_valid_out[20] [0]),
    .B(net1200),
    .Y(_2508_));
 sg13g2_nor2_1 _4159_ (.A(_2505_),
    .B(_2508_),
    .Y(_2509_));
 sg13g2_o21ai_1 _4160_ (.B1(_2457_),
    .Y(_2510_),
    .A1(\s0.was_valid_out[20] [0]),
    .A2(net1207));
 sg13g2_o21ai_1 _4161_ (.B1(_2510_),
    .Y(_2511_),
    .A1(net1195),
    .A2(_2503_));
 sg13g2_nor2_1 _4162_ (.A(_2509_),
    .B(_2511_),
    .Y(_2512_));
 sg13g2_o21ai_1 _4163_ (.B1(net1291),
    .Y(_2513_),
    .A1(net372),
    .A2(_2507_));
 sg13g2_nor2_1 _4164_ (.A(_2512_),
    .B(_2513_),
    .Y(_0001_));
 sg13g2_nor2_1 _4165_ (.A(net1217),
    .B(_2507_),
    .Y(_0002_));
 sg13g2_nor2b_1 _4166_ (.A(net1190),
    .B_N(net1073),
    .Y(_2514_));
 sg13g2_and2_1 _4167_ (.A(net1190),
    .B(\s0.data_out[20][0] ),
    .X(_2515_));
 sg13g2_o21ai_1 _4168_ (.B1(net1202),
    .Y(_2516_),
    .A1(_2514_),
    .A2(_2515_));
 sg13g2_nor2b_1 _4169_ (.A(net368),
    .B_N(net1206),
    .Y(_2517_));
 sg13g2_nor2_1 _4170_ (.A(net1206),
    .B(\s0.data_out[20][0] ),
    .Y(_2518_));
 sg13g2_nor3_1 _4171_ (.A(net1202),
    .B(_2517_),
    .C(_2518_),
    .Y(_2519_));
 sg13g2_nor2_1 _4172_ (.A(net1216),
    .B(_2519_),
    .Y(_2520_));
 sg13g2_a22oi_1 _4173_ (.Y(_0003_),
    .B1(_2516_),
    .B2(_2520_),
    .A2(_2482_),
    .A1(net1216));
 sg13g2_and2_1 _4174_ (.A(net1190),
    .B(\s0.data_out[20][1] ),
    .X(_2521_));
 sg13g2_nor2b_1 _4175_ (.A(net1190),
    .B_N(net1069),
    .Y(_2522_));
 sg13g2_o21ai_1 _4176_ (.B1(net1202),
    .Y(_2523_),
    .A1(_2521_),
    .A2(_2522_));
 sg13g2_a21oi_1 _4177_ (.A1(net1206),
    .A2(_2481_),
    .Y(_2524_),
    .B1(net1202));
 sg13g2_o21ai_1 _4178_ (.B1(_2524_),
    .Y(_2525_),
    .A1(net1206),
    .A2(\s0.data_out[20][1] ));
 sg13g2_nand3_1 _4179_ (.B(_2523_),
    .C(_2525_),
    .A(net1285),
    .Y(_2526_));
 sg13g2_o21ai_1 _4180_ (.B1(_2526_),
    .Y(_2527_),
    .A1(net1285),
    .A2(net370));
 sg13g2_inv_1 _4181_ (.Y(_0004_),
    .A(net371));
 sg13g2_and2_1 _4182_ (.A(net1191),
    .B(\s0.data_out[20][2] ),
    .X(_2528_));
 sg13g2_nor2b_1 _4183_ (.A(net1191),
    .B_N(net1065),
    .Y(_2529_));
 sg13g2_o21ai_1 _4184_ (.B1(net1202),
    .Y(_2530_),
    .A1(_2528_),
    .A2(_2529_));
 sg13g2_a21oi_1 _4185_ (.A1(net1206),
    .A2(_2479_),
    .Y(_2531_),
    .B1(net1203));
 sg13g2_o21ai_1 _4186_ (.B1(_2531_),
    .Y(_2532_),
    .A1(net1206),
    .A2(\s0.data_out[20][2] ));
 sg13g2_nand3_1 _4187_ (.B(_2530_),
    .C(_2532_),
    .A(net1285),
    .Y(_2533_));
 sg13g2_o21ai_1 _4188_ (.B1(_2533_),
    .Y(_2534_),
    .A1(net1285),
    .A2(net388));
 sg13g2_inv_1 _4189_ (.Y(_0005_),
    .A(net389));
 sg13g2_and2_1 _4190_ (.A(net1190),
    .B(\s0.data_out[20][3] ),
    .X(_2535_));
 sg13g2_nor2b_1 _4191_ (.A(net1190),
    .B_N(net1061),
    .Y(_2536_));
 sg13g2_o21ai_1 _4192_ (.B1(net1202),
    .Y(_2537_),
    .A1(_2535_),
    .A2(_2536_));
 sg13g2_nor2b_1 _4193_ (.A(net366),
    .B_N(net1206),
    .Y(_2538_));
 sg13g2_nor2_1 _4194_ (.A(net1206),
    .B(\s0.data_out[20][3] ),
    .Y(_2539_));
 sg13g2_nor3_1 _4195_ (.A(net1202),
    .B(_2538_),
    .C(_2539_),
    .Y(_2540_));
 sg13g2_nor2_1 _4196_ (.A(net1216),
    .B(_2540_),
    .Y(_2541_));
 sg13g2_a22oi_1 _4197_ (.Y(_0006_),
    .B1(_2537_),
    .B2(_2541_),
    .A2(_2478_),
    .A1(net1216));
 sg13g2_and2_1 _4198_ (.A(net1196),
    .B(\s0.data_out[20][4] ),
    .X(_2542_));
 sg13g2_nor2b_1 _4199_ (.A(net1195),
    .B_N(net1057),
    .Y(_2543_));
 sg13g2_o21ai_1 _4200_ (.B1(net1204),
    .Y(_2544_),
    .A1(_2542_),
    .A2(_2543_));
 sg13g2_nor2b_1 _4201_ (.A(net359),
    .B_N(net1207),
    .Y(_2545_));
 sg13g2_nor2_1 _4202_ (.A(net1207),
    .B(\s0.data_out[20][4] ),
    .Y(_2546_));
 sg13g2_nor3_1 _4203_ (.A(net1205),
    .B(_2545_),
    .C(_2546_),
    .Y(_2547_));
 sg13g2_nor2_1 _4204_ (.A(net1217),
    .B(_2547_),
    .Y(_2548_));
 sg13g2_a22oi_1 _4205_ (.Y(_0007_),
    .B1(_2544_),
    .B2(_2548_),
    .A2(_2477_),
    .A1(net1217));
 sg13g2_and2_1 _4206_ (.A(net1196),
    .B(\s0.data_out[20][5] ),
    .X(_2549_));
 sg13g2_nor2b_1 _4207_ (.A(net1195),
    .B_N(net1053),
    .Y(_2550_));
 sg13g2_o21ai_1 _4208_ (.B1(net1205),
    .Y(_2551_),
    .A1(_2549_),
    .A2(_2550_));
 sg13g2_nor2b_1 _4209_ (.A(net361),
    .B_N(\s0.valid_out[21] [0]),
    .Y(_2552_));
 sg13g2_nor2_1 _4210_ (.A(\s0.valid_out[21] [0]),
    .B(\s0.data_out[20][5] ),
    .Y(_2553_));
 sg13g2_nor3_1 _4211_ (.A(net1204),
    .B(_2552_),
    .C(_2553_),
    .Y(_2554_));
 sg13g2_nor2_1 _4212_ (.A(net1217),
    .B(_2554_),
    .Y(_2555_));
 sg13g2_a22oi_1 _4213_ (.Y(_0008_),
    .B1(_2551_),
    .B2(_2555_),
    .A2(_2475_),
    .A1(net1217));
 sg13g2_and2_1 _4214_ (.A(net1195),
    .B(\s0.data_out[20][6] ),
    .X(_2556_));
 sg13g2_nor2b_1 _4215_ (.A(net1195),
    .B_N(net1049),
    .Y(_2557_));
 sg13g2_o21ai_1 _4216_ (.B1(net1204),
    .Y(_2558_),
    .A1(_2556_),
    .A2(_2557_));
 sg13g2_nor2b_1 _4217_ (.A(net356),
    .B_N(net1207),
    .Y(_2559_));
 sg13g2_nor2_1 _4218_ (.A(\s0.valid_out[21] [0]),
    .B(\s0.data_out[20][6] ),
    .Y(_2560_));
 sg13g2_nor3_1 _4219_ (.A(net1204),
    .B(_2559_),
    .C(_2560_),
    .Y(_2561_));
 sg13g2_nor2_1 _4220_ (.A(net1216),
    .B(_2561_),
    .Y(_2562_));
 sg13g2_a22oi_1 _4221_ (.Y(_0009_),
    .B1(_2558_),
    .B2(_2562_),
    .A2(_2473_),
    .A1(net1216));
 sg13g2_and2_1 _4222_ (.A(net1192),
    .B(\s0.data_out[20][7] ),
    .X(_2563_));
 sg13g2_nor2b_1 _4223_ (.A(net1192),
    .B_N(net1045),
    .Y(_2564_));
 sg13g2_o21ai_1 _4224_ (.B1(net1203),
    .Y(_2565_),
    .A1(_2563_),
    .A2(_2564_));
 sg13g2_nor2b_1 _4225_ (.A(net364),
    .B_N(net1207),
    .Y(_2566_));
 sg13g2_nor2_1 _4226_ (.A(net1207),
    .B(\s0.data_out[20][7] ),
    .Y(_2567_));
 sg13g2_nor3_1 _4227_ (.A(net1203),
    .B(_2566_),
    .C(_2567_),
    .Y(_2568_));
 sg13g2_nor2_1 _4228_ (.A(net1216),
    .B(_2568_),
    .Y(_2569_));
 sg13g2_a22oi_1 _4229_ (.Y(_0010_),
    .B1(_2565_),
    .B2(_2569_),
    .A2(_2472_),
    .A1(net1216));
 sg13g2_nand2_1 _4230_ (.Y(_2570_),
    .A(net1198),
    .B(net490));
 sg13g2_o21ai_1 _4231_ (.B1(_2570_),
    .Y(_2571_),
    .A1(net1198),
    .A2(_2479_));
 sg13g2_a21oi_1 _4232_ (.A1(net1191),
    .A2(_2571_),
    .Y(_2572_),
    .B1(_2529_));
 sg13g2_o21ai_1 _4233_ (.B1(_2532_),
    .Y(_2573_),
    .A1(_2457_),
    .A2(_2572_));
 sg13g2_mux2_1 _4234_ (.A0(\s0.data_out[21][1] ),
    .A1(\s0.data_out[20][1] ),
    .S(net1198),
    .X(_2574_));
 sg13g2_a21oi_1 _4235_ (.A1(net1190),
    .A2(_2574_),
    .Y(_2575_),
    .B1(_2522_));
 sg13g2_nand2b_1 _4236_ (.Y(_2576_),
    .B(net1203),
    .A_N(_2575_));
 sg13g2_nand3_1 _4237_ (.B(_2525_),
    .C(_2576_),
    .A(net1273),
    .Y(_2577_));
 sg13g2_mux2_1 _4238_ (.A0(\s0.data_out[21][0] ),
    .A1(\s0.data_out[20][0] ),
    .S(net1198),
    .X(_2578_));
 sg13g2_a21o_1 _4239_ (.A2(_2578_),
    .A1(net1190),
    .B1(_2514_),
    .X(_2579_));
 sg13g2_a21oi_1 _4240_ (.A1(net1202),
    .A2(_2579_),
    .Y(_2580_),
    .B1(_2519_));
 sg13g2_nor2_1 _4241_ (.A(net1281),
    .B(_2580_),
    .Y(_2581_));
 sg13g2_a21oi_1 _4242_ (.A1(_2525_),
    .A2(_2576_),
    .Y(_2582_),
    .B1(net1273));
 sg13g2_a221oi_1 _4243_ (.B2(_2581_),
    .C1(_2582_),
    .B1(_2577_),
    .A1(net1211),
    .Y(_2583_),
    .A2(_2573_));
 sg13g2_nand2_1 _4244_ (.Y(_2584_),
    .A(net1198),
    .B(net560));
 sg13g2_mux2_1 _4245_ (.A0(\s0.data_out[21][3] ),
    .A1(\s0.data_out[20][3] ),
    .S(net1198),
    .X(_2585_));
 sg13g2_a21o_1 _4246_ (.A2(_2585_),
    .A1(net1191),
    .B1(_2536_),
    .X(_2586_));
 sg13g2_a21oi_1 _4247_ (.A1(net1203),
    .A2(_2586_),
    .Y(_2587_),
    .B1(_2540_));
 sg13g2_nand2_1 _4248_ (.Y(_2588_),
    .A(net1260),
    .B(_2587_));
 sg13g2_o21ai_1 _4249_ (.B1(_2588_),
    .Y(_2589_),
    .A1(net1211),
    .A2(_2573_));
 sg13g2_nor2_1 _4250_ (.A(_2583_),
    .B(_2589_),
    .Y(_2590_));
 sg13g2_nand2_1 _4251_ (.Y(_2591_),
    .A(net1198),
    .B(net523));
 sg13g2_mux2_1 _4252_ (.A0(\s0.data_out[21][7] ),
    .A1(\s0.data_out[20][7] ),
    .S(net1198),
    .X(_2592_));
 sg13g2_a21o_1 _4253_ (.A2(_2592_),
    .A1(net1192),
    .B1(_2564_),
    .X(_2593_));
 sg13g2_a21oi_1 _4254_ (.A1(net1203),
    .A2(_2593_),
    .Y(_2594_),
    .B1(_2568_));
 sg13g2_nand2_1 _4255_ (.Y(_2595_),
    .A(net1200),
    .B(net592));
 sg13g2_mux2_1 _4256_ (.A0(\s0.data_out[21][6] ),
    .A1(\s0.data_out[20][6] ),
    .S(net1200),
    .X(_2596_));
 sg13g2_a21o_1 _4257_ (.A2(_2596_),
    .A1(net1195),
    .B1(_2557_),
    .X(_2597_));
 sg13g2_a21oi_1 _4258_ (.A1(net1204),
    .A2(_2597_),
    .Y(_2598_),
    .B1(_2561_));
 sg13g2_a22oi_1 _4259_ (.Y(_2599_),
    .B1(_2598_),
    .B2(net1239),
    .A2(_2594_),
    .A1(net1231));
 sg13g2_nor2_1 _4260_ (.A(net1231),
    .B(_2594_),
    .Y(_2600_));
 sg13g2_or2_1 _4261_ (.X(_2601_),
    .B(_2598_),
    .A(net1239));
 sg13g2_nand3b_1 _4262_ (.B(_2601_),
    .C(_2599_),
    .Y(_2602_),
    .A_N(_2600_));
 sg13g2_mux2_1 _4263_ (.A0(\s0.data_out[21][4] ),
    .A1(\s0.data_out[20][4] ),
    .S(net1200),
    .X(_2603_));
 sg13g2_a21o_1 _4264_ (.A2(_2603_),
    .A1(net1195),
    .B1(_2543_),
    .X(_2604_));
 sg13g2_a21oi_1 _4265_ (.A1(net1204),
    .A2(_2604_),
    .Y(_2605_),
    .B1(_2547_));
 sg13g2_nand2_1 _4266_ (.Y(_2606_),
    .A(net1254),
    .B(_2605_));
 sg13g2_mux2_1 _4267_ (.A0(\s0.data_out[21][5] ),
    .A1(\s0.data_out[20][5] ),
    .S(net1200),
    .X(_2607_));
 sg13g2_a21o_1 _4268_ (.A2(_2607_),
    .A1(net1196),
    .B1(_2550_),
    .X(_2608_));
 sg13g2_a21oi_1 _4269_ (.A1(net1205),
    .A2(_2608_),
    .Y(_2609_),
    .B1(_2554_));
 sg13g2_nand2_1 _4270_ (.Y(_2610_),
    .A(net1246),
    .B(_2609_));
 sg13g2_nand2_1 _4271_ (.Y(_2611_),
    .A(_2606_),
    .B(_2610_));
 sg13g2_nor2_1 _4272_ (.A(net1260),
    .B(_2587_),
    .Y(_2612_));
 sg13g2_nor2_1 _4273_ (.A(net1246),
    .B(_2609_),
    .Y(_2613_));
 sg13g2_nor2_1 _4274_ (.A(_2612_),
    .B(_2613_),
    .Y(_2614_));
 sg13g2_o21ai_1 _4275_ (.B1(_2614_),
    .Y(_2615_),
    .A1(net1254),
    .A2(_2605_));
 sg13g2_or4_1 _4276_ (.A(_2590_),
    .B(_2602_),
    .C(_2611_),
    .D(_2615_),
    .X(_2616_));
 sg13g2_nor2_1 _4277_ (.A(_2599_),
    .B(_2600_),
    .Y(_2617_));
 sg13g2_o21ai_1 _4278_ (.B1(_2610_),
    .Y(_2618_),
    .A1(_2606_),
    .A2(_2613_));
 sg13g2_nor2b_1 _4279_ (.A(_2602_),
    .B_N(_2618_),
    .Y(_2619_));
 sg13g2_nor3_1 _4280_ (.A(_2507_),
    .B(_2617_),
    .C(_2619_),
    .Y(_2620_));
 sg13g2_nand2_1 _4281_ (.Y(_2621_),
    .A(net1223),
    .B(net1292));
 sg13g2_or2_1 _4282_ (.X(_2622_),
    .B(net1208),
    .A(net306));
 sg13g2_a21oi_1 _4283_ (.A1(_2616_),
    .A2(_2620_),
    .Y(_0011_),
    .B1(_2622_));
 sg13g2_and2_1 _4284_ (.A(net1285),
    .B(net301),
    .X(_0012_));
 sg13g2_o21ai_1 _4285_ (.B1(net1196),
    .Y(_2623_),
    .A1(net1225),
    .A2(net1182));
 sg13g2_nand2_1 _4286_ (.Y(_2624_),
    .A(net1222),
    .B(net1189));
 sg13g2_nand2b_1 _4287_ (.Y(_2625_),
    .B(_2624_),
    .A_N(_2623_));
 sg13g2_o21ai_1 _4288_ (.B1(_2625_),
    .Y(_2626_),
    .A1(net1197),
    .A2(_2504_));
 sg13g2_nor2_1 _4289_ (.A(net323),
    .B(net1188),
    .Y(_2627_));
 sg13g2_or2_1 _4290_ (.X(_2628_),
    .B(_2627_),
    .A(_2625_));
 sg13g2_nor2_1 _4291_ (.A(net1182),
    .B(_2623_),
    .Y(_2629_));
 sg13g2_o21ai_1 _4292_ (.B1(_2456_),
    .Y(_2630_),
    .A1(net323),
    .A2(net1201));
 sg13g2_nor2b_1 _4293_ (.A(_2629_),
    .B_N(_2630_),
    .Y(_2631_));
 sg13g2_o21ai_1 _4294_ (.B1(net1289),
    .Y(_2632_),
    .A1(net435),
    .A2(_2626_));
 sg13g2_a21oi_1 _4295_ (.A1(_2628_),
    .A2(_2631_),
    .Y(_0013_),
    .B1(_2632_));
 sg13g2_nor2_1 _4296_ (.A(net1217),
    .B(_2626_),
    .Y(_0014_));
 sg13g2_mux2_1 _4297_ (.A0(\s0.data_out[19][0] ),
    .A1(\s0.data_out[20][0] ),
    .S(net1199),
    .X(_2633_));
 sg13g2_nand2_1 _4298_ (.Y(_2634_),
    .A(net931),
    .B(_2633_));
 sg13g2_and2_1 _4299_ (.A(net1178),
    .B(\s0.data_out[19][0] ),
    .X(_2635_));
 sg13g2_nor2b_1 _4300_ (.A(net1178),
    .B_N(net1073),
    .Y(_2636_));
 sg13g2_o21ai_1 _4301_ (.B1(net1193),
    .Y(_2637_),
    .A1(_2635_),
    .A2(_2636_));
 sg13g2_nand3_1 _4302_ (.B(_2634_),
    .C(_2637_),
    .A(net1286),
    .Y(_2638_));
 sg13g2_o21ai_1 _4303_ (.B1(_2638_),
    .Y(_2639_),
    .A1(net1285),
    .A2(net462));
 sg13g2_inv_1 _4304_ (.Y(_0015_),
    .A(_2639_));
 sg13g2_mux2_1 _4305_ (.A0(\s0.data_out[19][1] ),
    .A1(\s0.data_out[20][1] ),
    .S(net1199),
    .X(_2640_));
 sg13g2_nand2_1 _4306_ (.Y(_2641_),
    .A(net931),
    .B(_2640_));
 sg13g2_and2_1 _4307_ (.A(net1178),
    .B(\s0.data_out[19][1] ),
    .X(_2642_));
 sg13g2_nor2b_1 _4308_ (.A(net1178),
    .B_N(net1069),
    .Y(_2643_));
 sg13g2_o21ai_1 _4309_ (.B1(net1193),
    .Y(_2644_),
    .A1(_2642_),
    .A2(_2643_));
 sg13g2_nand3_1 _4310_ (.B(_2641_),
    .C(_2644_),
    .A(net1286),
    .Y(_2645_));
 sg13g2_o21ai_1 _4311_ (.B1(_2645_),
    .Y(_2646_),
    .A1(net1286),
    .A2(net455));
 sg13g2_inv_1 _4312_ (.Y(_0016_),
    .A(_2646_));
 sg13g2_nand2b_1 _4313_ (.Y(_2647_),
    .B(net475),
    .A_N(net1199));
 sg13g2_a21oi_1 _4314_ (.A1(_2570_),
    .A2(_2647_),
    .Y(_2648_),
    .B1(net1193));
 sg13g2_nor2b_1 _4315_ (.A(net1178),
    .B_N(net1065),
    .Y(_2649_));
 sg13g2_a21oi_1 _4316_ (.A1(net1179),
    .A2(net475),
    .Y(_2650_),
    .B1(_2649_));
 sg13g2_o21ai_1 _4317_ (.B1(net1286),
    .Y(_2651_),
    .A1(net931),
    .A2(_2650_));
 sg13g2_or2_1 _4318_ (.X(_2652_),
    .B(net490),
    .A(net1285));
 sg13g2_o21ai_1 _4319_ (.B1(_2652_),
    .Y(_2653_),
    .A1(_2648_),
    .A2(_2651_));
 sg13g2_inv_1 _4320_ (.Y(_0017_),
    .A(_2653_));
 sg13g2_nand2b_1 _4321_ (.Y(_2654_),
    .B(\s0.data_out[19][3] ),
    .A_N(net1199));
 sg13g2_a21oi_1 _4322_ (.A1(_2584_),
    .A2(_2654_),
    .Y(_2655_),
    .B1(net1193));
 sg13g2_nor2b_1 _4323_ (.A(net1179),
    .B_N(net1061),
    .Y(_2656_));
 sg13g2_a21oi_1 _4324_ (.A1(net1179),
    .A2(\s0.data_out[19][3] ),
    .Y(_2657_),
    .B1(_2656_));
 sg13g2_o21ai_1 _4325_ (.B1(net1286),
    .Y(_2658_),
    .A1(net931),
    .A2(_2657_));
 sg13g2_or2_1 _4326_ (.X(_2659_),
    .B(net560),
    .A(net1286));
 sg13g2_o21ai_1 _4327_ (.B1(_2659_),
    .Y(_2660_),
    .A1(_2655_),
    .A2(_2658_));
 sg13g2_inv_1 _4328_ (.Y(_0018_),
    .A(net561));
 sg13g2_mux2_1 _4329_ (.A0(\s0.data_out[19][4] ),
    .A1(\s0.data_out[20][4] ),
    .S(net1200),
    .X(_2661_));
 sg13g2_nand2_1 _4330_ (.Y(_2662_),
    .A(net931),
    .B(_2661_));
 sg13g2_and2_1 _4331_ (.A(net1182),
    .B(\s0.data_out[19][4] ),
    .X(_2663_));
 sg13g2_nor2b_1 _4332_ (.A(net1182),
    .B_N(net1057),
    .Y(_2664_));
 sg13g2_o21ai_1 _4333_ (.B1(net1196),
    .Y(_2665_),
    .A1(_2663_),
    .A2(_2664_));
 sg13g2_nand3_1 _4334_ (.B(_2662_),
    .C(_2665_),
    .A(net1289),
    .Y(_2666_));
 sg13g2_o21ai_1 _4335_ (.B1(_2666_),
    .Y(_2667_),
    .A1(net1289),
    .A2(net469));
 sg13g2_inv_1 _4336_ (.Y(_0019_),
    .A(_2667_));
 sg13g2_mux2_1 _4337_ (.A0(\s0.data_out[19][5] ),
    .A1(\s0.data_out[20][5] ),
    .S(net1200),
    .X(_2668_));
 sg13g2_nand2_1 _4338_ (.Y(_2669_),
    .A(net931),
    .B(_2668_));
 sg13g2_and2_1 _4339_ (.A(net1183),
    .B(\s0.data_out[19][5] ),
    .X(_2670_));
 sg13g2_nor2b_1 _4340_ (.A(net1182),
    .B_N(net1053),
    .Y(_2671_));
 sg13g2_o21ai_1 _4341_ (.B1(net1196),
    .Y(_2672_),
    .A1(_2670_),
    .A2(_2671_));
 sg13g2_nand3_1 _4342_ (.B(_2669_),
    .C(_2672_),
    .A(net1289),
    .Y(_2673_));
 sg13g2_o21ai_1 _4343_ (.B1(_2673_),
    .Y(_2674_),
    .A1(net1285),
    .A2(net395));
 sg13g2_inv_1 _4344_ (.Y(_0020_),
    .A(_2674_));
 sg13g2_nand2b_1 _4345_ (.Y(_2675_),
    .B(net551),
    .A_N(net1201));
 sg13g2_a21oi_1 _4346_ (.A1(_2595_),
    .A2(_2675_),
    .Y(_2676_),
    .B1(net1197));
 sg13g2_nor2b_1 _4347_ (.A(net1182),
    .B_N(net1049),
    .Y(_2677_));
 sg13g2_a21oi_1 _4348_ (.A1(net1182),
    .A2(net551),
    .Y(_2678_),
    .B1(_2677_));
 sg13g2_o21ai_1 _4349_ (.B1(net1286),
    .Y(_2679_),
    .A1(_2456_),
    .A2(_2678_));
 sg13g2_or2_1 _4350_ (.X(_2680_),
    .B(net592),
    .A(net1288));
 sg13g2_o21ai_1 _4351_ (.B1(_2680_),
    .Y(_2681_),
    .A1(_2676_),
    .A2(_2679_));
 sg13g2_inv_1 _4352_ (.Y(_0021_),
    .A(_2681_));
 sg13g2_nand2b_1 _4353_ (.Y(_2682_),
    .B(\s0.data_out[19][7] ),
    .A_N(net1199));
 sg13g2_a21oi_1 _4354_ (.A1(_2591_),
    .A2(_2682_),
    .Y(_2683_),
    .B1(net1194));
 sg13g2_nor2b_1 _4355_ (.A(net1180),
    .B_N(net1045),
    .Y(_2684_));
 sg13g2_a21oi_1 _4356_ (.A1(net1180),
    .A2(\s0.data_out[19][7] ),
    .Y(_2685_),
    .B1(_2684_));
 sg13g2_o21ai_1 _4357_ (.B1(net1286),
    .Y(_2686_),
    .A1(net931),
    .A2(_2685_));
 sg13g2_or2_1 _4358_ (.X(_2687_),
    .B(net523),
    .A(net1288));
 sg13g2_o21ai_1 _4359_ (.B1(_2687_),
    .Y(_2688_),
    .A1(_2683_),
    .A2(_2686_));
 sg13g2_inv_1 _4360_ (.Y(_0022_),
    .A(net524));
 sg13g2_mux2_1 _4361_ (.A0(\s0.data_out[20][2] ),
    .A1(\s0.data_out[19][2] ),
    .S(net1186),
    .X(_2689_));
 sg13g2_a21o_1 _4362_ (.A2(_2689_),
    .A1(net1178),
    .B1(_2649_),
    .X(_2690_));
 sg13g2_a21oi_1 _4363_ (.A1(net1193),
    .A2(_2690_),
    .Y(_2691_),
    .B1(_2648_));
 sg13g2_or2_1 _4364_ (.X(_2692_),
    .B(_2691_),
    .A(net1268));
 sg13g2_nand2_1 _4365_ (.Y(_2693_),
    .A(net1187),
    .B(\s0.data_out[19][1] ));
 sg13g2_mux2_1 _4366_ (.A0(\s0.data_out[20][1] ),
    .A1(\s0.data_out[19][1] ),
    .S(net1186),
    .X(_2694_));
 sg13g2_a21oi_1 _4367_ (.A1(net1178),
    .A2(_2694_),
    .Y(_2695_),
    .B1(_2643_));
 sg13g2_nand2b_1 _4368_ (.Y(_2696_),
    .B(net1193),
    .A_N(_2695_));
 sg13g2_and2_1 _4369_ (.A(_2641_),
    .B(_2696_),
    .X(_2697_));
 sg13g2_mux2_1 _4370_ (.A0(\s0.data_out[20][0] ),
    .A1(\s0.data_out[19][0] ),
    .S(net1186),
    .X(_2698_));
 sg13g2_a21oi_1 _4371_ (.A1(net1178),
    .A2(_2698_),
    .Y(_2699_),
    .B1(_2636_));
 sg13g2_nand2b_1 _4372_ (.Y(_2700_),
    .B(net1193),
    .A_N(_2699_));
 sg13g2_a221oi_1 _4373_ (.B2(_2634_),
    .C1(net1281),
    .B1(_2700_),
    .A1(net1273),
    .Y(_2701_),
    .A2(_2697_));
 sg13g2_o21ai_1 _4374_ (.B1(_2692_),
    .Y(_2702_),
    .A1(net1273),
    .A2(_2697_));
 sg13g2_nand2_1 _4375_ (.Y(_2703_),
    .A(net1186),
    .B(net567));
 sg13g2_mux2_1 _4376_ (.A0(\s0.data_out[20][3] ),
    .A1(\s0.data_out[19][3] ),
    .S(net1186),
    .X(_2704_));
 sg13g2_a21o_1 _4377_ (.A2(_2704_),
    .A1(net1179),
    .B1(_2656_),
    .X(_2705_));
 sg13g2_a21oi_1 _4378_ (.A1(net1193),
    .A2(_2705_),
    .Y(_2706_),
    .B1(_2655_));
 sg13g2_a22oi_1 _4379_ (.Y(_2707_),
    .B1(_2706_),
    .B2(net1260),
    .A2(_2691_),
    .A1(net1268));
 sg13g2_o21ai_1 _4380_ (.B1(_2707_),
    .Y(_2708_),
    .A1(_2701_),
    .A2(_2702_));
 sg13g2_nand2_1 _4381_ (.Y(_2709_),
    .A(net1186),
    .B(net574));
 sg13g2_mux2_1 _4382_ (.A0(\s0.data_out[20][7] ),
    .A1(\s0.data_out[19][7] ),
    .S(net1186),
    .X(_2710_));
 sg13g2_a21o_1 _4383_ (.A2(_2710_),
    .A1(net1180),
    .B1(_2684_),
    .X(_2711_));
 sg13g2_a21oi_1 _4384_ (.A1(net1197),
    .A2(_2711_),
    .Y(_2712_),
    .B1(_2683_));
 sg13g2_nand2_1 _4385_ (.Y(_2713_),
    .A(net1188),
    .B(net551));
 sg13g2_mux2_1 _4386_ (.A0(\s0.data_out[20][6] ),
    .A1(\s0.data_out[19][6] ),
    .S(net1188),
    .X(_2714_));
 sg13g2_a21o_1 _4387_ (.A2(_2714_),
    .A1(net1182),
    .B1(_2677_),
    .X(_2715_));
 sg13g2_a21oi_1 _4388_ (.A1(net1197),
    .A2(_2715_),
    .Y(_2716_),
    .B1(_2676_));
 sg13g2_a22oi_1 _4389_ (.Y(_2717_),
    .B1(_2716_),
    .B2(net1239),
    .A2(_2712_),
    .A1(net1231));
 sg13g2_or2_1 _4390_ (.X(_2718_),
    .B(_2712_),
    .A(net1231));
 sg13g2_or2_1 _4391_ (.X(_2719_),
    .B(_2716_),
    .A(net1239));
 sg13g2_and3_1 _4392_ (.X(_2720_),
    .A(_2717_),
    .B(_2718_),
    .C(_2719_));
 sg13g2_mux2_1 _4393_ (.A0(\s0.data_out[20][4] ),
    .A1(\s0.data_out[19][4] ),
    .S(net1188),
    .X(_2721_));
 sg13g2_a21oi_1 _4394_ (.A1(net1183),
    .A2(_2721_),
    .Y(_2722_),
    .B1(_2664_));
 sg13g2_o21ai_1 _4395_ (.B1(_2662_),
    .Y(_2723_),
    .A1(net931),
    .A2(_2722_));
 sg13g2_nand2_1 _4396_ (.Y(_2724_),
    .A(net1188),
    .B(net586));
 sg13g2_mux2_1 _4397_ (.A0(\s0.data_out[20][5] ),
    .A1(\s0.data_out[19][5] ),
    .S(net1188),
    .X(_2725_));
 sg13g2_a21oi_1 _4398_ (.A1(net1183),
    .A2(_2725_),
    .Y(_2726_),
    .B1(_2671_));
 sg13g2_nand2b_1 _4399_ (.Y(_2727_),
    .B(net1196),
    .A_N(_2726_));
 sg13g2_nand3_1 _4400_ (.B(_2669_),
    .C(_2727_),
    .A(net1246),
    .Y(_2728_));
 sg13g2_a21oi_1 _4401_ (.A1(_2669_),
    .A2(_2727_),
    .Y(_2729_),
    .B1(net1246));
 sg13g2_nor2_1 _4402_ (.A(net1260),
    .B(_2706_),
    .Y(_2730_));
 sg13g2_nor2_1 _4403_ (.A(_2729_),
    .B(_2730_),
    .Y(_2731_));
 sg13g2_xnor2_1 _4404_ (.Y(_2732_),
    .A(net1254),
    .B(_2723_));
 sg13g2_and4_1 _4405_ (.A(_2720_),
    .B(_2728_),
    .C(_2731_),
    .D(_2732_),
    .X(_2733_));
 sg13g2_or3_1 _4406_ (.A(net1214),
    .B(_2723_),
    .C(_2729_),
    .X(_2734_));
 sg13g2_nand2_1 _4407_ (.Y(_2735_),
    .A(_2728_),
    .B(_2734_));
 sg13g2_nand2b_1 _4408_ (.Y(_2736_),
    .B(_2718_),
    .A_N(_2717_));
 sg13g2_a221oi_1 _4409_ (.B2(_2720_),
    .C1(_2626_),
    .B1(_2735_),
    .A1(_2708_),
    .Y(_2737_),
    .A2(_2733_));
 sg13g2_or2_1 _4410_ (.X(_2738_),
    .B(net1208),
    .A(net301));
 sg13g2_a21oi_1 _4411_ (.A1(_2736_),
    .A2(_2737_),
    .Y(_0023_),
    .B1(_2738_));
 sg13g2_and2_1 _4412_ (.A(net1295),
    .B(net297),
    .X(_0024_));
 sg13g2_o21ai_1 _4413_ (.B1(net1183),
    .Y(_2739_),
    .A1(net1226),
    .A2(net1170));
 sg13g2_nor2b_1 _4414_ (.A(net1226),
    .B_N(net1176),
    .Y(_2740_));
 sg13g2_nor2_1 _4415_ (.A(_2739_),
    .B(_2740_),
    .Y(_2741_));
 sg13g2_a21oi_1 _4416_ (.A1(net926),
    .A2(_2624_),
    .Y(_2742_),
    .B1(_2741_));
 sg13g2_o21ai_1 _4417_ (.B1(_2741_),
    .Y(_2743_),
    .A1(\s0.was_valid_out[18] [0]),
    .A2(net1176));
 sg13g2_nor2_1 _4418_ (.A(net1172),
    .B(_2739_),
    .Y(_2744_));
 sg13g2_o21ai_1 _4419_ (.B1(net927),
    .Y(_2745_),
    .A1(\s0.was_valid_out[18] [0]),
    .A2(net1188));
 sg13g2_nand2_1 _4420_ (.Y(_2746_),
    .A(_2743_),
    .B(_2745_));
 sg13g2_o21ai_1 _4421_ (.B1(net1290),
    .Y(_2747_),
    .A1(_2744_),
    .A2(_2746_));
 sg13g2_a21oi_1 _4422_ (.A1(_2447_),
    .A2(_2742_),
    .Y(_0025_),
    .B1(_2747_));
 sg13g2_and2_1 _4423_ (.A(net1290),
    .B(_2742_),
    .X(_0026_));
 sg13g2_mux2_1 _4424_ (.A0(\s0.data_out[18][0] ),
    .A1(\s0.data_out[19][0] ),
    .S(net1187),
    .X(_2748_));
 sg13g2_nand2_1 _4425_ (.Y(_2749_),
    .A(net926),
    .B(_2748_));
 sg13g2_and2_1 _4426_ (.A(net1167),
    .B(\s0.data_out[18][0] ),
    .X(_2750_));
 sg13g2_nor2b_1 _4427_ (.A(net1167),
    .B_N(net1073),
    .Y(_2751_));
 sg13g2_o21ai_1 _4428_ (.B1(net1181),
    .Y(_2752_),
    .A1(_2750_),
    .A2(_2751_));
 sg13g2_nand3_1 _4429_ (.B(_2749_),
    .C(_2752_),
    .A(net1287),
    .Y(_2753_));
 sg13g2_o21ai_1 _4430_ (.B1(_2753_),
    .Y(_2754_),
    .A1(net1287),
    .A2(net410));
 sg13g2_inv_1 _4431_ (.Y(_0027_),
    .A(_2754_));
 sg13g2_o21ai_1 _4432_ (.B1(_2693_),
    .Y(_2755_),
    .A1(net1187),
    .A2(_2484_));
 sg13g2_nand2_1 _4433_ (.Y(_2756_),
    .A(net926),
    .B(_2755_));
 sg13g2_nor2_1 _4434_ (.A(net925),
    .B(_2484_),
    .Y(_2757_));
 sg13g2_nor2b_1 _4435_ (.A(net1167),
    .B_N(net1069),
    .Y(_2758_));
 sg13g2_o21ai_1 _4436_ (.B1(net1181),
    .Y(_2759_),
    .A1(_2757_),
    .A2(_2758_));
 sg13g2_nand3_1 _4437_ (.B(_2756_),
    .C(_2759_),
    .A(net1302),
    .Y(_2760_));
 sg13g2_o21ai_1 _4438_ (.B1(_2760_),
    .Y(_2761_),
    .A1(net1287),
    .A2(net464));
 sg13g2_inv_1 _4439_ (.Y(_0028_),
    .A(_2761_));
 sg13g2_mux2_1 _4440_ (.A0(\s0.data_out[18][2] ),
    .A1(\s0.data_out[19][2] ),
    .S(net1186),
    .X(_2762_));
 sg13g2_nand2_1 _4441_ (.Y(_2763_),
    .A(net926),
    .B(_2762_));
 sg13g2_and2_1 _4442_ (.A(net1167),
    .B(\s0.data_out[18][2] ),
    .X(_2764_));
 sg13g2_nor2b_1 _4443_ (.A(net1168),
    .B_N(net1065),
    .Y(_2765_));
 sg13g2_o21ai_1 _4444_ (.B1(net1181),
    .Y(_2766_),
    .A1(_2764_),
    .A2(_2765_));
 sg13g2_nand3_1 _4445_ (.B(_2763_),
    .C(_2766_),
    .A(net1287),
    .Y(_2767_));
 sg13g2_o21ai_1 _4446_ (.B1(_2767_),
    .Y(_2768_),
    .A1(net1287),
    .A2(net475));
 sg13g2_inv_1 _4447_ (.Y(_0029_),
    .A(_2768_));
 sg13g2_nand2b_1 _4448_ (.Y(_2769_),
    .B(net478),
    .A_N(net1187));
 sg13g2_a21oi_1 _4449_ (.A1(_2703_),
    .A2(_2769_),
    .Y(_2770_),
    .B1(net1181));
 sg13g2_nor2b_1 _4450_ (.A(net1167),
    .B_N(net1061),
    .Y(_2771_));
 sg13g2_a21oi_1 _4451_ (.A1(net1167),
    .A2(net478),
    .Y(_2772_),
    .B1(_2771_));
 sg13g2_o21ai_1 _4452_ (.B1(net1287),
    .Y(_2773_),
    .A1(net926),
    .A2(_2772_));
 sg13g2_or2_1 _4453_ (.X(_2774_),
    .B(net567),
    .A(net1287));
 sg13g2_o21ai_1 _4454_ (.B1(_2774_),
    .Y(_2775_),
    .A1(_2770_),
    .A2(_2773_));
 sg13g2_inv_1 _4455_ (.Y(_0030_),
    .A(_2775_));
 sg13g2_mux2_1 _4456_ (.A0(\s0.data_out[18][4] ),
    .A1(\s0.data_out[19][4] ),
    .S(net1188),
    .X(_2776_));
 sg13g2_nand2_1 _4457_ (.Y(_2777_),
    .A(net927),
    .B(_2776_));
 sg13g2_and2_1 _4458_ (.A(net1170),
    .B(\s0.data_out[18][4] ),
    .X(_2778_));
 sg13g2_nor2b_1 _4459_ (.A(net1170),
    .B_N(net1057),
    .Y(_2779_));
 sg13g2_o21ai_1 _4460_ (.B1(net1183),
    .Y(_2780_),
    .A1(_2778_),
    .A2(_2779_));
 sg13g2_nand3_1 _4461_ (.B(_2777_),
    .C(_2780_),
    .A(net1289),
    .Y(_2781_));
 sg13g2_o21ai_1 _4462_ (.B1(_2781_),
    .Y(_2782_),
    .A1(net1289),
    .A2(net414));
 sg13g2_inv_1 _4463_ (.Y(_0031_),
    .A(_2782_));
 sg13g2_nand2b_1 _4464_ (.Y(_2783_),
    .B(net570),
    .A_N(net1189));
 sg13g2_a21oi_1 _4465_ (.A1(_2724_),
    .A2(_2783_),
    .Y(_2784_),
    .B1(net1184));
 sg13g2_nor2b_1 _4466_ (.A(net1170),
    .B_N(net1053),
    .Y(_2785_));
 sg13g2_a21oi_1 _4467_ (.A1(net1172),
    .A2(net570),
    .Y(_2786_),
    .B1(_2785_));
 sg13g2_o21ai_1 _4468_ (.B1(net1289),
    .Y(_2787_),
    .A1(net927),
    .A2(_2786_));
 sg13g2_or2_1 _4469_ (.X(_2788_),
    .B(net586),
    .A(net1290));
 sg13g2_o21ai_1 _4470_ (.B1(_2788_),
    .Y(_2789_),
    .A1(_2784_),
    .A2(_2787_));
 sg13g2_inv_1 _4471_ (.Y(_0032_),
    .A(_2789_));
 sg13g2_nand2b_1 _4472_ (.Y(_2790_),
    .B(\s0.data_out[18][6] ),
    .A_N(net1189));
 sg13g2_a21oi_1 _4473_ (.A1(_2713_),
    .A2(_2790_),
    .Y(_2791_),
    .B1(net1184));
 sg13g2_nor2b_1 _4474_ (.A(net1170),
    .B_N(net1049),
    .Y(_2792_));
 sg13g2_a21oi_1 _4475_ (.A1(net1170),
    .A2(\s0.data_out[18][6] ),
    .Y(_2793_),
    .B1(_2792_));
 sg13g2_o21ai_1 _4476_ (.B1(net1287),
    .Y(_2794_),
    .A1(net927),
    .A2(_2793_));
 sg13g2_or2_1 _4477_ (.X(_2795_),
    .B(net551),
    .A(net1288));
 sg13g2_o21ai_1 _4478_ (.B1(_2795_),
    .Y(_2796_),
    .A1(_2791_),
    .A2(_2794_));
 sg13g2_inv_1 _4479_ (.Y(_0033_),
    .A(net552));
 sg13g2_nand2b_1 _4480_ (.Y(_2797_),
    .B(\s0.data_out[18][7] ),
    .A_N(net1187));
 sg13g2_a21oi_1 _4481_ (.A1(_2709_),
    .A2(_2797_),
    .Y(_2798_),
    .B1(net1185));
 sg13g2_nor2b_1 _4482_ (.A(net1168),
    .B_N(net1045),
    .Y(_2799_));
 sg13g2_a21oi_1 _4483_ (.A1(net1168),
    .A2(\s0.data_out[18][7] ),
    .Y(_2800_),
    .B1(_2799_));
 sg13g2_o21ai_1 _4484_ (.B1(net1288),
    .Y(_2801_),
    .A1(net926),
    .A2(_2800_));
 sg13g2_or2_1 _4485_ (.X(_2802_),
    .B(net574),
    .A(net1288));
 sg13g2_o21ai_1 _4486_ (.B1(_2802_),
    .Y(_2803_),
    .A1(_2798_),
    .A2(_2801_));
 sg13g2_inv_1 _4487_ (.Y(_0034_),
    .A(net575));
 sg13g2_nand2_1 _4488_ (.Y(_2804_),
    .A(net1174),
    .B(net498));
 sg13g2_o21ai_1 _4489_ (.B1(_2804_),
    .Y(_2805_),
    .A1(net1174),
    .A2(_2483_));
 sg13g2_a21oi_1 _4490_ (.A1(net1168),
    .A2(_2805_),
    .Y(_2806_),
    .B1(_2765_));
 sg13g2_o21ai_1 _4491_ (.B1(_2763_),
    .Y(_2807_),
    .A1(net926),
    .A2(_2806_));
 sg13g2_nand2_1 _4492_ (.Y(_2808_),
    .A(net1174),
    .B(net493));
 sg13g2_mux2_1 _4493_ (.A0(\s0.data_out[19][1] ),
    .A1(\s0.data_out[18][1] ),
    .S(net1174),
    .X(_2809_));
 sg13g2_a21oi_1 _4494_ (.A1(net1168),
    .A2(_2809_),
    .Y(_2810_),
    .B1(_2758_));
 sg13g2_nand2b_1 _4495_ (.Y(_2811_),
    .B(net1181),
    .A_N(_2810_));
 sg13g2_nand3_1 _4496_ (.B(_2756_),
    .C(_2811_),
    .A(net1275),
    .Y(_2812_));
 sg13g2_a21oi_1 _4497_ (.A1(_2756_),
    .A2(_2811_),
    .Y(_2813_),
    .B1(net1275));
 sg13g2_mux2_1 _4498_ (.A0(\s0.data_out[19][0] ),
    .A1(\s0.data_out[18][0] ),
    .S(net1174),
    .X(_2814_));
 sg13g2_a21oi_1 _4499_ (.A1(net1167),
    .A2(_2814_),
    .Y(_2815_),
    .B1(_2751_));
 sg13g2_o21ai_1 _4500_ (.B1(_2749_),
    .Y(_2816_),
    .A1(net926),
    .A2(_2815_));
 sg13g2_nor2b_1 _4501_ (.A(net1284),
    .B_N(_2816_),
    .Y(_2817_));
 sg13g2_a221oi_1 _4502_ (.B2(_2817_),
    .C1(_2813_),
    .B1(_2812_),
    .A1(net1212),
    .Y(_2818_),
    .A2(_2807_));
 sg13g2_mux2_1 _4503_ (.A0(\s0.data_out[19][3] ),
    .A1(\s0.data_out[18][3] ),
    .S(net1174),
    .X(_2819_));
 sg13g2_a21o_1 _4504_ (.A2(_2819_),
    .A1(net1167),
    .B1(_2771_),
    .X(_2820_));
 sg13g2_a21oi_1 _4505_ (.A1(net1181),
    .A2(_2820_),
    .Y(_2821_),
    .B1(_2770_));
 sg13g2_nand2_1 _4506_ (.Y(_2822_),
    .A(net1262),
    .B(_2821_));
 sg13g2_o21ai_1 _4507_ (.B1(_2822_),
    .Y(_2823_),
    .A1(net1212),
    .A2(_2807_));
 sg13g2_nor2_1 _4508_ (.A(_2818_),
    .B(_2823_),
    .Y(_2824_));
 sg13g2_nand2_1 _4509_ (.Y(_2825_),
    .A(net1174),
    .B(net579));
 sg13g2_mux2_1 _4510_ (.A0(\s0.data_out[19][7] ),
    .A1(\s0.data_out[18][7] ),
    .S(net1174),
    .X(_2826_));
 sg13g2_a21o_1 _4511_ (.A2(_2826_),
    .A1(net1168),
    .B1(_2799_),
    .X(_2827_));
 sg13g2_a21oi_1 _4512_ (.A1(net1183),
    .A2(_2827_),
    .Y(_2828_),
    .B1(_2798_));
 sg13g2_nand2_1 _4513_ (.Y(_2829_),
    .A(net1176),
    .B(net558));
 sg13g2_mux2_1 _4514_ (.A0(\s0.data_out[19][6] ),
    .A1(\s0.data_out[18][6] ),
    .S(net1176),
    .X(_2830_));
 sg13g2_a21o_1 _4515_ (.A2(_2830_),
    .A1(net1170),
    .B1(_2792_),
    .X(_2831_));
 sg13g2_a21oi_1 _4516_ (.A1(net1184),
    .A2(_2831_),
    .Y(_2832_),
    .B1(_2791_));
 sg13g2_a22oi_1 _4517_ (.Y(_2833_),
    .B1(_2832_),
    .B2(net1240),
    .A2(_2828_),
    .A1(net1231));
 sg13g2_nor2_1 _4518_ (.A(net1239),
    .B(_2832_),
    .Y(_2834_));
 sg13g2_or2_1 _4519_ (.X(_0272_),
    .B(_2828_),
    .A(net1231));
 sg13g2_nand3b_1 _4520_ (.B(_0272_),
    .C(_2833_),
    .Y(_0273_),
    .A_N(_2834_));
 sg13g2_nand2_1 _4521_ (.Y(_0274_),
    .A(net1176),
    .B(net570));
 sg13g2_mux2_1 _4522_ (.A0(\s0.data_out[19][5] ),
    .A1(\s0.data_out[18][5] ),
    .S(net1176),
    .X(_0275_));
 sg13g2_a21o_1 _4523_ (.A2(_0275_),
    .A1(net1172),
    .B1(_2785_),
    .X(_0276_));
 sg13g2_a21oi_1 _4524_ (.A1(net1184),
    .A2(_0276_),
    .Y(_0277_),
    .B1(_2784_));
 sg13g2_nand2_1 _4525_ (.Y(_0278_),
    .A(net1248),
    .B(_0277_));
 sg13g2_mux2_1 _4526_ (.A0(\s0.data_out[19][4] ),
    .A1(\s0.data_out[18][4] ),
    .S(net1176),
    .X(_0279_));
 sg13g2_a21oi_1 _4527_ (.A1(net1170),
    .A2(_0279_),
    .Y(_0280_),
    .B1(_2779_));
 sg13g2_nand2b_1 _4528_ (.Y(_0281_),
    .B(net1183),
    .A_N(_0280_));
 sg13g2_nand3_1 _4529_ (.B(_2777_),
    .C(_0281_),
    .A(net1254),
    .Y(_0282_));
 sg13g2_a21oi_1 _4530_ (.A1(_2777_),
    .A2(_0281_),
    .Y(_0283_),
    .B1(net1254));
 sg13g2_nor2_1 _4531_ (.A(net1248),
    .B(_0277_),
    .Y(_0284_));
 sg13g2_nor2_1 _4532_ (.A(net1262),
    .B(_2821_),
    .Y(_0285_));
 sg13g2_nor3_1 _4533_ (.A(_0283_),
    .B(_0284_),
    .C(_0285_),
    .Y(_0286_));
 sg13g2_nand3_1 _4534_ (.B(_0282_),
    .C(_0286_),
    .A(_0278_),
    .Y(_0287_));
 sg13g2_or3_1 _4535_ (.A(_2824_),
    .B(_0273_),
    .C(_0287_),
    .X(_0288_));
 sg13g2_o21ai_1 _4536_ (.B1(_0278_),
    .Y(_0289_),
    .A1(_0282_),
    .A2(_0284_));
 sg13g2_nand2b_1 _4537_ (.Y(_0290_),
    .B(_0289_),
    .A_N(_0273_));
 sg13g2_nand2b_1 _4538_ (.Y(_0291_),
    .B(_0272_),
    .A_N(_2833_));
 sg13g2_and3_1 _4539_ (.X(_0292_),
    .A(_2742_),
    .B(_0290_),
    .C(_0291_));
 sg13g2_or2_1 _4540_ (.X(_0293_),
    .B(net1208),
    .A(net305));
 sg13g2_a21oi_1 _4541_ (.A1(_0288_),
    .A2(_0292_),
    .Y(_0035_),
    .B1(_0293_));
 sg13g2_and2_1 _4542_ (.A(net1303),
    .B(net304),
    .X(_0036_));
 sg13g2_o21ai_1 _4543_ (.B1(net1171),
    .Y(_0294_),
    .A1(net1226),
    .A2(net1158));
 sg13g2_nor2b_1 _4544_ (.A(net1226),
    .B_N(net1163),
    .Y(_0295_));
 sg13g2_nor2_1 _4545_ (.A(_0294_),
    .B(_0295_),
    .Y(_0296_));
 sg13g2_inv_1 _4546_ (.Y(_0297_),
    .A(_0296_));
 sg13g2_o21ai_1 _4547_ (.B1(_0297_),
    .Y(_0298_),
    .A1(net1171),
    .A2(_2740_));
 sg13g2_or2_1 _4548_ (.X(_0299_),
    .B(net1166),
    .A(net375));
 sg13g2_o21ai_1 _4549_ (.B1(net925),
    .Y(_0300_),
    .A1(net375),
    .A2(net1177));
 sg13g2_o21ai_1 _4550_ (.B1(_0300_),
    .Y(_0301_),
    .A1(net1158),
    .A2(_0294_));
 sg13g2_a21oi_1 _4551_ (.A1(_0296_),
    .A2(_0299_),
    .Y(_0302_),
    .B1(_0301_));
 sg13g2_o21ai_1 _4552_ (.B1(net1303),
    .Y(_0303_),
    .A1(net406),
    .A2(_0298_));
 sg13g2_nor2_1 _4553_ (.A(_0302_),
    .B(_0303_),
    .Y(_0037_));
 sg13g2_nor2_1 _4554_ (.A(net1219),
    .B(_0298_),
    .Y(_0038_));
 sg13g2_mux2_1 _4555_ (.A0(\s0.data_out[17][0] ),
    .A1(\s0.data_out[18][0] ),
    .S(net1175),
    .X(_0304_));
 sg13g2_nand2_1 _4556_ (.Y(_0305_),
    .A(net925),
    .B(_0304_));
 sg13g2_and2_1 _4557_ (.A(net1155),
    .B(\s0.data_out[17][0] ),
    .X(_0306_));
 sg13g2_nor2b_1 _4558_ (.A(net1155),
    .B_N(net1076),
    .Y(_0307_));
 sg13g2_o21ai_1 _4559_ (.B1(net1169),
    .Y(_0308_),
    .A1(_0306_),
    .A2(_0307_));
 sg13g2_nand3_1 _4560_ (.B(_0305_),
    .C(_0308_),
    .A(net1301),
    .Y(_0309_));
 sg13g2_o21ai_1 _4561_ (.B1(_0309_),
    .Y(_0310_),
    .A1(net1301),
    .A2(net460));
 sg13g2_inv_1 _4562_ (.Y(_0039_),
    .A(_0310_));
 sg13g2_nand2b_1 _4563_ (.Y(_0311_),
    .B(\s0.data_out[17][1] ),
    .A_N(net1175));
 sg13g2_a21oi_1 _4564_ (.A1(_2808_),
    .A2(_0311_),
    .Y(_0312_),
    .B1(net1169));
 sg13g2_nor2b_1 _4565_ (.A(net1155),
    .B_N(net1072),
    .Y(_0313_));
 sg13g2_a21oi_1 _4566_ (.A1(net1156),
    .A2(\s0.data_out[17][1] ),
    .Y(_0314_),
    .B1(_0313_));
 sg13g2_o21ai_1 _4567_ (.B1(net1301),
    .Y(_0315_),
    .A1(net925),
    .A2(_0314_));
 sg13g2_nand2_1 _4568_ (.Y(_0316_),
    .A(net1219),
    .B(_2484_));
 sg13g2_o21ai_1 _4569_ (.B1(_0316_),
    .Y(_0317_),
    .A1(_0312_),
    .A2(_0315_));
 sg13g2_inv_1 _4570_ (.Y(_0040_),
    .A(net494));
 sg13g2_nand2b_1 _4571_ (.Y(_0318_),
    .B(\s0.data_out[17][2] ),
    .A_N(net1175));
 sg13g2_a21oi_1 _4572_ (.A1(_2804_),
    .A2(_0318_),
    .Y(_0319_),
    .B1(net1169));
 sg13g2_nor2b_1 _4573_ (.A(net1155),
    .B_N(net1068),
    .Y(_0320_));
 sg13g2_a21oi_1 _4574_ (.A1(net1155),
    .A2(\s0.data_out[17][2] ),
    .Y(_0321_),
    .B1(_0320_));
 sg13g2_o21ai_1 _4575_ (.B1(net1301),
    .Y(_0322_),
    .A1(net925),
    .A2(_0321_));
 sg13g2_or2_1 _4576_ (.X(_0323_),
    .B(net498),
    .A(net1302));
 sg13g2_o21ai_1 _4577_ (.B1(_0323_),
    .Y(_0324_),
    .A1(_0319_),
    .A2(_0322_));
 sg13g2_inv_1 _4578_ (.Y(_0041_),
    .A(net499));
 sg13g2_mux2_1 _4579_ (.A0(\s0.data_out[17][3] ),
    .A1(\s0.data_out[18][3] ),
    .S(net1175),
    .X(_0325_));
 sg13g2_nand2_1 _4580_ (.Y(_0326_),
    .A(net925),
    .B(_0325_));
 sg13g2_and2_1 _4581_ (.A(net1156),
    .B(\s0.data_out[17][3] ),
    .X(_0327_));
 sg13g2_nor2b_1 _4582_ (.A(net1156),
    .B_N(net1061),
    .Y(_0328_));
 sg13g2_o21ai_1 _4583_ (.B1(net1169),
    .Y(_0329_),
    .A1(_0327_),
    .A2(_0328_));
 sg13g2_nand3_1 _4584_ (.B(_0326_),
    .C(_0329_),
    .A(net1301),
    .Y(_0330_));
 sg13g2_o21ai_1 _4585_ (.B1(_0330_),
    .Y(_0331_),
    .A1(net1301),
    .A2(net478));
 sg13g2_inv_1 _4586_ (.Y(_0042_),
    .A(_0331_));
 sg13g2_mux2_1 _4587_ (.A0(\s0.data_out[17][4] ),
    .A1(\s0.data_out[18][4] ),
    .S(net1176),
    .X(_0332_));
 sg13g2_nand2_1 _4588_ (.Y(_0333_),
    .A(net925),
    .B(_0332_));
 sg13g2_and2_1 _4589_ (.A(net1158),
    .B(\s0.data_out[17][4] ),
    .X(_0334_));
 sg13g2_nor2b_1 _4590_ (.A(net1158),
    .B_N(net1058),
    .Y(_0335_));
 sg13g2_o21ai_1 _4591_ (.B1(net1171),
    .Y(_0336_),
    .A1(_0334_),
    .A2(_0335_));
 sg13g2_nand3_1 _4592_ (.B(_0333_),
    .C(_0336_),
    .A(net1303),
    .Y(_0337_));
 sg13g2_o21ai_1 _4593_ (.B1(_0337_),
    .Y(_0338_),
    .A1(net1303),
    .A2(net325));
 sg13g2_inv_1 _4594_ (.Y(_0043_),
    .A(_0338_));
 sg13g2_nand2b_1 _4595_ (.Y(_0339_),
    .B(\s0.data_out[17][5] ),
    .A_N(net1177));
 sg13g2_a21oi_1 _4596_ (.A1(_0274_),
    .A2(_0339_),
    .Y(_0340_),
    .B1(net1172));
 sg13g2_nor2b_1 _4597_ (.A(net1159),
    .B_N(net1054),
    .Y(_0341_));
 sg13g2_a21oi_1 _4598_ (.A1(net1159),
    .A2(\s0.data_out[17][5] ),
    .Y(_0342_),
    .B1(_0341_));
 sg13g2_o21ai_1 _4599_ (.B1(net1303),
    .Y(_0343_),
    .A1(_2461_),
    .A2(_0342_));
 sg13g2_or2_1 _4600_ (.X(_0344_),
    .B(net570),
    .A(net1303));
 sg13g2_o21ai_1 _4601_ (.B1(_0344_),
    .Y(_0345_),
    .A1(_0340_),
    .A2(_0343_));
 sg13g2_inv_1 _4602_ (.Y(_0044_),
    .A(net571));
 sg13g2_nand2b_1 _4603_ (.Y(_0346_),
    .B(\s0.data_out[17][6] ),
    .A_N(net1177));
 sg13g2_a21oi_1 _4604_ (.A1(_2829_),
    .A2(_0346_),
    .Y(_0347_),
    .B1(net1171));
 sg13g2_nor2b_1 _4605_ (.A(net1158),
    .B_N(net1050),
    .Y(_0348_));
 sg13g2_a21oi_1 _4606_ (.A1(net1158),
    .A2(\s0.data_out[17][6] ),
    .Y(_0349_),
    .B1(_0348_));
 sg13g2_o21ai_1 _4607_ (.B1(net1301),
    .Y(_0350_),
    .A1(_2461_),
    .A2(_0349_));
 sg13g2_or2_1 _4608_ (.X(_0351_),
    .B(net558),
    .A(net1302));
 sg13g2_o21ai_1 _4609_ (.B1(_0351_),
    .Y(_0352_),
    .A1(_0347_),
    .A2(_0350_));
 sg13g2_inv_1 _4610_ (.Y(_0045_),
    .A(net559));
 sg13g2_nand2b_1 _4611_ (.Y(_0353_),
    .B(net341),
    .A_N(net1175));
 sg13g2_a21oi_1 _4612_ (.A1(_2825_),
    .A2(_0353_),
    .Y(_0354_),
    .B1(net1173));
 sg13g2_nor2b_1 _4613_ (.A(net1157),
    .B_N(net1046),
    .Y(_0355_));
 sg13g2_a21oi_1 _4614_ (.A1(net1157),
    .A2(net341),
    .Y(_0356_),
    .B1(_0355_));
 sg13g2_o21ai_1 _4615_ (.B1(net1301),
    .Y(_0357_),
    .A1(net925),
    .A2(_0356_));
 sg13g2_or2_1 _4616_ (.X(_0358_),
    .B(net579),
    .A(net1302));
 sg13g2_o21ai_1 _4617_ (.B1(_0358_),
    .Y(_0359_),
    .A1(_0354_),
    .A2(_0357_));
 sg13g2_inv_1 _4618_ (.Y(_0046_),
    .A(net580));
 sg13g2_nand2_1 _4619_ (.Y(_0360_),
    .A(net1164),
    .B(net530));
 sg13g2_mux2_1 _4620_ (.A0(\s0.data_out[18][2] ),
    .A1(\s0.data_out[17][2] ),
    .S(net1163),
    .X(_0361_));
 sg13g2_a21o_1 _4621_ (.A2(_0361_),
    .A1(net1155),
    .B1(_0320_),
    .X(_0362_));
 sg13g2_a21oi_1 _4622_ (.A1(net1169),
    .A2(_0362_),
    .Y(_0363_),
    .B1(_0319_));
 sg13g2_or2_1 _4623_ (.X(_0364_),
    .B(_0363_),
    .A(net1269));
 sg13g2_nand2_1 _4624_ (.Y(_0365_),
    .A(net1163),
    .B(net496));
 sg13g2_o21ai_1 _4625_ (.B1(_0365_),
    .Y(_0366_),
    .A1(net1163),
    .A2(_2484_));
 sg13g2_a21o_1 _4626_ (.A2(_0366_),
    .A1(net1156),
    .B1(_0313_),
    .X(_0367_));
 sg13g2_a21oi_1 _4627_ (.A1(net1169),
    .A2(_0367_),
    .Y(_0368_),
    .B1(_0312_));
 sg13g2_mux2_1 _4628_ (.A0(\s0.data_out[18][0] ),
    .A1(\s0.data_out[17][0] ),
    .S(net1163),
    .X(_0369_));
 sg13g2_a21oi_1 _4629_ (.A1(net1155),
    .A2(_0369_),
    .Y(_0370_),
    .B1(_0307_));
 sg13g2_nand2b_1 _4630_ (.Y(_0371_),
    .B(net1169),
    .A_N(_0370_));
 sg13g2_o21ai_1 _4631_ (.B1(_0364_),
    .Y(_0372_),
    .A1(net1275),
    .A2(_0368_));
 sg13g2_a221oi_1 _4632_ (.B2(_0305_),
    .C1(net1281),
    .B1(_0371_),
    .A1(net1275),
    .Y(_0373_),
    .A2(_0368_));
 sg13g2_nand2_1 _4633_ (.Y(_0374_),
    .A(net1164),
    .B(\s0.data_out[17][3] ));
 sg13g2_mux2_1 _4634_ (.A0(\s0.data_out[18][3] ),
    .A1(\s0.data_out[17][3] ),
    .S(net1163),
    .X(_0375_));
 sg13g2_a21oi_1 _4635_ (.A1(net1155),
    .A2(_0375_),
    .Y(_0376_),
    .B1(_0328_));
 sg13g2_nand2b_1 _4636_ (.Y(_0377_),
    .B(net1169),
    .A_N(_0376_));
 sg13g2_and2_1 _4637_ (.A(_0326_),
    .B(_0377_),
    .X(_0378_));
 sg13g2_a22oi_1 _4638_ (.Y(_0379_),
    .B1(_0378_),
    .B2(net1262),
    .A2(_0363_),
    .A1(net1269));
 sg13g2_o21ai_1 _4639_ (.B1(_0379_),
    .Y(_0380_),
    .A1(_0372_),
    .A2(_0373_));
 sg13g2_nand2_1 _4640_ (.Y(_0381_),
    .A(net1164),
    .B(net341));
 sg13g2_mux2_1 _4641_ (.A0(\s0.data_out[18][7] ),
    .A1(\s0.data_out[17][7] ),
    .S(net1163),
    .X(_0382_));
 sg13g2_a21o_1 _4642_ (.A2(_0382_),
    .A1(net1157),
    .B1(_0355_),
    .X(_0383_));
 sg13g2_a21oi_1 _4643_ (.A1(net1171),
    .A2(_0383_),
    .Y(_0384_),
    .B1(_0354_));
 sg13g2_nand2_1 _4644_ (.Y(_0385_),
    .A(net1165),
    .B(net572));
 sg13g2_mux2_1 _4645_ (.A0(\s0.data_out[18][6] ),
    .A1(\s0.data_out[17][6] ),
    .S(net1166),
    .X(_0386_));
 sg13g2_a21o_1 _4646_ (.A2(_0386_),
    .A1(net1158),
    .B1(_0348_),
    .X(_0387_));
 sg13g2_a21oi_1 _4647_ (.A1(net1171),
    .A2(_0387_),
    .Y(_0388_),
    .B1(_0347_));
 sg13g2_a22oi_1 _4648_ (.Y(_0389_),
    .B1(_0388_),
    .B2(net1240),
    .A2(_0384_),
    .A1(net1233));
 sg13g2_nor2_1 _4649_ (.A(net1240),
    .B(_0388_),
    .Y(_0390_));
 sg13g2_or2_1 _4650_ (.X(_0391_),
    .B(_0384_),
    .A(net1233));
 sg13g2_nand3b_1 _4651_ (.B(_0391_),
    .C(_0389_),
    .Y(_0392_),
    .A_N(_0390_));
 sg13g2_nand2_1 _4652_ (.Y(_0393_),
    .A(net1165),
    .B(net582));
 sg13g2_mux2_1 _4653_ (.A0(\s0.data_out[18][5] ),
    .A1(\s0.data_out[17][5] ),
    .S(net1166),
    .X(_0394_));
 sg13g2_a21o_1 _4654_ (.A2(_0394_),
    .A1(net1159),
    .B1(_0341_),
    .X(_0395_));
 sg13g2_a21oi_1 _4655_ (.A1(net1172),
    .A2(_0395_),
    .Y(_0396_),
    .B1(_0340_));
 sg13g2_nand2_1 _4656_ (.Y(_0397_),
    .A(net1248),
    .B(_0396_));
 sg13g2_o21ai_1 _4657_ (.B1(_0397_),
    .Y(_0398_),
    .A1(net1262),
    .A2(_0378_));
 sg13g2_mux2_1 _4658_ (.A0(\s0.data_out[18][4] ),
    .A1(\s0.data_out[17][4] ),
    .S(net1163),
    .X(_0399_));
 sg13g2_a21oi_1 _4659_ (.A1(net1158),
    .A2(_0399_),
    .Y(_0400_),
    .B1(_0335_));
 sg13g2_nand2b_1 _4660_ (.Y(_0401_),
    .B(net1171),
    .A_N(_0400_));
 sg13g2_a21o_1 _4661_ (.A2(_0401_),
    .A1(_0333_),
    .B1(net1255),
    .X(_0402_));
 sg13g2_nand3_1 _4662_ (.B(_0333_),
    .C(_0401_),
    .A(net1255),
    .Y(_0403_));
 sg13g2_nor2_1 _4663_ (.A(net1248),
    .B(_0396_),
    .Y(_0404_));
 sg13g2_nor3_1 _4664_ (.A(_0392_),
    .B(_0398_),
    .C(_0404_),
    .Y(_0405_));
 sg13g2_nand4_1 _4665_ (.B(_0402_),
    .C(_0403_),
    .A(_0380_),
    .Y(_0406_),
    .D(_0405_));
 sg13g2_o21ai_1 _4666_ (.B1(_0397_),
    .Y(_0407_),
    .A1(_0403_),
    .A2(_0404_));
 sg13g2_nor2b_1 _4667_ (.A(_0392_),
    .B_N(_0407_),
    .Y(_0408_));
 sg13g2_nor2b_1 _4668_ (.A(_0389_),
    .B_N(_0391_),
    .Y(_0409_));
 sg13g2_nor3_1 _4669_ (.A(_0298_),
    .B(_0408_),
    .C(_0409_),
    .Y(_0410_));
 sg13g2_or2_1 _4670_ (.X(_0411_),
    .B(net1210),
    .A(net304));
 sg13g2_a21oi_1 _4671_ (.A1(_0406_),
    .A2(_0410_),
    .Y(_0047_),
    .B1(_0411_));
 sg13g2_and2_1 _4672_ (.A(net1306),
    .B(net308),
    .X(_0048_));
 sg13g2_o21ai_1 _4673_ (.B1(net1161),
    .Y(_0412_),
    .A1(net1226),
    .A2(net1146));
 sg13g2_a21oi_1 _4674_ (.A1(net1222),
    .A2(net1151),
    .Y(_0413_),
    .B1(_0412_));
 sg13g2_inv_1 _4675_ (.Y(_0414_),
    .A(_0413_));
 sg13g2_o21ai_1 _4676_ (.B1(_0413_),
    .Y(_0415_),
    .A1(net321),
    .A2(net1151));
 sg13g2_nor2_1 _4677_ (.A(net1146),
    .B(_0412_),
    .Y(_0416_));
 sg13g2_o21ai_1 _4678_ (.B1(net924),
    .Y(_0417_),
    .A1(net321),
    .A2(net1165));
 sg13g2_nor2b_1 _4679_ (.A(_0416_),
    .B_N(_0417_),
    .Y(_0418_));
 sg13g2_o21ai_1 _4680_ (.B1(_0414_),
    .Y(_0419_),
    .A1(net1159),
    .A2(_0295_));
 sg13g2_o21ai_1 _4681_ (.B1(net1306),
    .Y(_0420_),
    .A1(net375),
    .A2(_0419_));
 sg13g2_a21oi_1 _4682_ (.A1(_0415_),
    .A2(_0418_),
    .Y(_0049_),
    .B1(_0420_));
 sg13g2_nor2_1 _4683_ (.A(net1219),
    .B(_0419_),
    .Y(_0050_));
 sg13g2_mux2_1 _4684_ (.A0(\s0.data_out[16][0] ),
    .A1(\s0.data_out[17][0] ),
    .S(net1164),
    .X(_0421_));
 sg13g2_nand2_1 _4685_ (.Y(_0422_),
    .A(net924),
    .B(_0421_));
 sg13g2_and2_1 _4686_ (.A(net1144),
    .B(\s0.data_out[16][0] ),
    .X(_0423_));
 sg13g2_nor2b_1 _4687_ (.A(net1144),
    .B_N(net1073),
    .Y(_0424_));
 sg13g2_o21ai_1 _4688_ (.B1(net1160),
    .Y(_0425_),
    .A1(_0423_),
    .A2(_0424_));
 sg13g2_nand3_1 _4689_ (.B(_0422_),
    .C(_0425_),
    .A(net1304),
    .Y(_0426_));
 sg13g2_o21ai_1 _4690_ (.B1(_0426_),
    .Y(_0427_),
    .A1(net1304),
    .A2(net468));
 sg13g2_inv_1 _4691_ (.Y(_0051_),
    .A(_0427_));
 sg13g2_nand2b_1 _4692_ (.Y(_0428_),
    .B(net476),
    .A_N(net1164));
 sg13g2_a21oi_1 _4693_ (.A1(_0365_),
    .A2(_0428_),
    .Y(_0429_),
    .B1(net1162));
 sg13g2_nor2b_1 _4694_ (.A(net1144),
    .B_N(net1069),
    .Y(_0430_));
 sg13g2_a21oi_1 _4695_ (.A1(net1144),
    .A2(net476),
    .Y(_0431_),
    .B1(_0430_));
 sg13g2_o21ai_1 _4696_ (.B1(net1304),
    .Y(_0432_),
    .A1(net924),
    .A2(_0431_));
 sg13g2_or2_1 _4697_ (.X(_0433_),
    .B(net496),
    .A(net1304));
 sg13g2_o21ai_1 _4698_ (.B1(_0433_),
    .Y(_0434_),
    .A1(_0429_),
    .A2(_0432_));
 sg13g2_inv_1 _4699_ (.Y(_0052_),
    .A(net497));
 sg13g2_nand2b_1 _4700_ (.Y(_0435_),
    .B(net422),
    .A_N(net1164));
 sg13g2_a21oi_1 _4701_ (.A1(_0360_),
    .A2(_0435_),
    .Y(_0436_),
    .B1(net1161));
 sg13g2_nor2b_1 _4702_ (.A(net1145),
    .B_N(net1065),
    .Y(_0437_));
 sg13g2_a21oi_1 _4703_ (.A1(net1144),
    .A2(net422),
    .Y(_0438_),
    .B1(_0437_));
 sg13g2_o21ai_1 _4704_ (.B1(net1304),
    .Y(_0439_),
    .A1(net924),
    .A2(_0438_));
 sg13g2_or2_1 _4705_ (.X(_0440_),
    .B(net530),
    .A(net1304));
 sg13g2_o21ai_1 _4706_ (.B1(_0440_),
    .Y(_0441_),
    .A1(_0436_),
    .A2(_0439_));
 sg13g2_inv_1 _4707_ (.Y(_0053_),
    .A(_0441_));
 sg13g2_o21ai_1 _4708_ (.B1(_0374_),
    .Y(_0442_),
    .A1(net1164),
    .A2(_2485_));
 sg13g2_nand2_1 _4709_ (.Y(_0443_),
    .A(net924),
    .B(_0442_));
 sg13g2_nor2_1 _4710_ (.A(net922),
    .B(_2485_),
    .Y(_0444_));
 sg13g2_nor2b_1 _4711_ (.A(net1147),
    .B_N(net1062),
    .Y(_0445_));
 sg13g2_o21ai_1 _4712_ (.B1(net1160),
    .Y(_0446_),
    .A1(_0444_),
    .A2(_0445_));
 sg13g2_nand3_1 _4713_ (.B(_0443_),
    .C(_0446_),
    .A(net1305),
    .Y(_0447_));
 sg13g2_o21ai_1 _4714_ (.B1(_0447_),
    .Y(_0448_),
    .A1(net1305),
    .A2(net480));
 sg13g2_inv_1 _4715_ (.Y(_0054_),
    .A(_0448_));
 sg13g2_mux2_1 _4716_ (.A0(\s0.data_out[16][4] ),
    .A1(\s0.data_out[17][4] ),
    .S(net1165),
    .X(_0449_));
 sg13g2_nand2_1 _4717_ (.Y(_0450_),
    .A(net924),
    .B(_0449_));
 sg13g2_and2_1 _4718_ (.A(net1146),
    .B(\s0.data_out[16][4] ),
    .X(_0451_));
 sg13g2_nor2b_1 _4719_ (.A(net1146),
    .B_N(net1057),
    .Y(_0452_));
 sg13g2_o21ai_1 _4720_ (.B1(net1161),
    .Y(_0453_),
    .A1(_0451_),
    .A2(_0452_));
 sg13g2_nand3_1 _4721_ (.B(_0450_),
    .C(_0453_),
    .A(net1306),
    .Y(_0454_));
 sg13g2_o21ai_1 _4722_ (.B1(_0454_),
    .Y(_0455_),
    .A1(net1306),
    .A2(net401));
 sg13g2_inv_1 _4723_ (.Y(_0055_),
    .A(_0455_));
 sg13g2_nand2b_1 _4724_ (.Y(_0456_),
    .B(net456),
    .A_N(net1165));
 sg13g2_a21oi_1 _4725_ (.A1(_0393_),
    .A2(_0456_),
    .Y(_0457_),
    .B1(net1162));
 sg13g2_nor2b_1 _4726_ (.A(net1146),
    .B_N(net1053),
    .Y(_0458_));
 sg13g2_a21oi_1 _4727_ (.A1(net1147),
    .A2(net456),
    .Y(_0459_),
    .B1(_0458_));
 sg13g2_o21ai_1 _4728_ (.B1(net1306),
    .Y(_0460_),
    .A1(_2462_),
    .A2(_0459_));
 sg13g2_or2_1 _4729_ (.X(_0461_),
    .B(net582),
    .A(net1306));
 sg13g2_o21ai_1 _4730_ (.B1(_0461_),
    .Y(_0462_),
    .A1(_0457_),
    .A2(_0460_));
 sg13g2_inv_1 _4731_ (.Y(_0056_),
    .A(net583));
 sg13g2_nand2b_1 _4732_ (.Y(_0463_),
    .B(net546),
    .A_N(net1165));
 sg13g2_a21oi_1 _4733_ (.A1(_0385_),
    .A2(_0463_),
    .Y(_0464_),
    .B1(net1161));
 sg13g2_nor2b_1 _4734_ (.A(net1147),
    .B_N(net1049),
    .Y(_0465_));
 sg13g2_a21oi_1 _4735_ (.A1(net1146),
    .A2(net546),
    .Y(_0466_),
    .B1(_0465_));
 sg13g2_o21ai_1 _4736_ (.B1(net1305),
    .Y(_0467_),
    .A1(_2462_),
    .A2(_0466_));
 sg13g2_or2_1 _4737_ (.X(_0468_),
    .B(net572),
    .A(net1304));
 sg13g2_o21ai_1 _4738_ (.B1(_0468_),
    .Y(_0469_),
    .A1(_0464_),
    .A2(_0467_));
 sg13g2_inv_1 _4739_ (.Y(_0057_),
    .A(_0469_));
 sg13g2_nand2b_1 _4740_ (.Y(_0470_),
    .B(\s0.data_out[16][7] ),
    .A_N(net1164));
 sg13g2_a21oi_1 _4741_ (.A1(_0381_),
    .A2(_0470_),
    .Y(_0471_),
    .B1(net1160));
 sg13g2_nor2b_1 _4742_ (.A(net1145),
    .B_N(net1045),
    .Y(_0472_));
 sg13g2_a21oi_1 _4743_ (.A1(net1145),
    .A2(net591),
    .Y(_0473_),
    .B1(_0472_));
 sg13g2_o21ai_1 _4744_ (.B1(net1304),
    .Y(_0474_),
    .A1(net924),
    .A2(_0473_));
 sg13g2_or2_1 _4745_ (.X(_0475_),
    .B(net341),
    .A(net1305));
 sg13g2_o21ai_1 _4746_ (.B1(_0475_),
    .Y(_0476_),
    .A1(net342),
    .A2(_0474_));
 sg13g2_inv_1 _4747_ (.Y(_0058_),
    .A(_0476_));
 sg13g2_mux2_1 _4748_ (.A0(\s0.data_out[17][2] ),
    .A1(\s0.data_out[16][2] ),
    .S(net1151),
    .X(_0477_));
 sg13g2_a21o_1 _4749_ (.A2(_0477_),
    .A1(net1144),
    .B1(_0437_),
    .X(_0478_));
 sg13g2_a21oi_1 _4750_ (.A1(net1160),
    .A2(_0478_),
    .Y(_0479_),
    .B1(_0436_));
 sg13g2_or2_1 _4751_ (.X(_0480_),
    .B(_0479_),
    .A(net1268));
 sg13g2_mux2_1 _4752_ (.A0(\s0.data_out[17][1] ),
    .A1(\s0.data_out[16][1] ),
    .S(net1151),
    .X(_0481_));
 sg13g2_a21o_1 _4753_ (.A2(_0481_),
    .A1(net1144),
    .B1(_0430_),
    .X(_0482_));
 sg13g2_a21oi_1 _4754_ (.A1(net1160),
    .A2(_0482_),
    .Y(_0483_),
    .B1(_0429_));
 sg13g2_mux2_1 _4755_ (.A0(\s0.data_out[17][0] ),
    .A1(\s0.data_out[16][0] ),
    .S(net1151),
    .X(_0484_));
 sg13g2_a21oi_1 _4756_ (.A1(net1144),
    .A2(_0484_),
    .Y(_0485_),
    .B1(_0424_));
 sg13g2_nand2b_1 _4757_ (.Y(_0486_),
    .B(net1160),
    .A_N(_0485_));
 sg13g2_a221oi_1 _4758_ (.B2(_0422_),
    .C1(net1282),
    .B1(_0486_),
    .A1(net1275),
    .Y(_0487_),
    .A2(_0483_));
 sg13g2_o21ai_1 _4759_ (.B1(_0480_),
    .Y(_0488_),
    .A1(net1277),
    .A2(_0483_));
 sg13g2_nand2_1 _4760_ (.Y(_0489_),
    .A(net1152),
    .B(net550));
 sg13g2_mux2_1 _4761_ (.A0(\s0.data_out[17][3] ),
    .A1(\s0.data_out[16][3] ),
    .S(net1151),
    .X(_0490_));
 sg13g2_a21oi_1 _4762_ (.A1(net1147),
    .A2(_0490_),
    .Y(_0491_),
    .B1(_0445_));
 sg13g2_nand2b_1 _4763_ (.Y(_0492_),
    .B(net1161),
    .A_N(_0491_));
 sg13g2_and2_1 _4764_ (.A(_0443_),
    .B(_0492_),
    .X(_0493_));
 sg13g2_a22oi_1 _4765_ (.Y(_0494_),
    .B1(_0493_),
    .B2(net1262),
    .A2(_0479_),
    .A1(net1268));
 sg13g2_o21ai_1 _4766_ (.B1(_0494_),
    .Y(_0495_),
    .A1(_0487_),
    .A2(_0488_));
 sg13g2_nand2_1 _4767_ (.Y(_0496_),
    .A(net1152),
    .B(net546));
 sg13g2_mux2_1 _4768_ (.A0(\s0.data_out[17][6] ),
    .A1(\s0.data_out[16][6] ),
    .S(net1154),
    .X(_0497_));
 sg13g2_a21o_1 _4769_ (.A2(_0497_),
    .A1(net1146),
    .B1(_0465_),
    .X(_0498_));
 sg13g2_a21oi_1 _4770_ (.A1(net1161),
    .A2(_0498_),
    .Y(_0499_),
    .B1(_0464_));
 sg13g2_nand2_1 _4771_ (.Y(_0500_),
    .A(net1152),
    .B(net591));
 sg13g2_mux2_1 _4772_ (.A0(\s0.data_out[17][7] ),
    .A1(\s0.data_out[16][7] ),
    .S(net1151),
    .X(_0501_));
 sg13g2_a21o_1 _4773_ (.A2(_0501_),
    .A1(net1145),
    .B1(_0472_),
    .X(_0502_));
 sg13g2_a21oi_1 _4774_ (.A1(net1160),
    .A2(_0502_),
    .Y(_0503_),
    .B1(_0471_));
 sg13g2_a22oi_1 _4775_ (.Y(_0504_),
    .B1(_0503_),
    .B2(net1233),
    .A2(_0499_),
    .A1(net1240));
 sg13g2_or2_1 _4776_ (.X(_0505_),
    .B(_0503_),
    .A(net1233));
 sg13g2_or2_1 _4777_ (.X(_0506_),
    .B(_0499_),
    .A(net1240));
 sg13g2_and3_1 _4778_ (.X(_0507_),
    .A(_0504_),
    .B(_0505_),
    .C(_0506_));
 sg13g2_nand3_1 _4779_ (.B(_0505_),
    .C(_0506_),
    .A(_0504_),
    .Y(_0508_));
 sg13g2_mux2_1 _4780_ (.A0(\s0.data_out[17][4] ),
    .A1(\s0.data_out[16][4] ),
    .S(net1151),
    .X(_0509_));
 sg13g2_a21oi_1 _4781_ (.A1(net1146),
    .A2(_0509_),
    .Y(_0510_),
    .B1(_0452_));
 sg13g2_o21ai_1 _4782_ (.B1(_0450_),
    .Y(_0511_),
    .A1(net924),
    .A2(_0510_));
 sg13g2_mux2_1 _4783_ (.A0(\s0.data_out[17][5] ),
    .A1(\s0.data_out[16][5] ),
    .S(net1154),
    .X(_0512_));
 sg13g2_a21o_1 _4784_ (.A2(_0512_),
    .A1(net1147),
    .B1(_0458_),
    .X(_0513_));
 sg13g2_a21oi_1 _4785_ (.A1(net1161),
    .A2(_0513_),
    .Y(_0514_),
    .B1(_0457_));
 sg13g2_nand2_1 _4786_ (.Y(_0515_),
    .A(net1248),
    .B(_0514_));
 sg13g2_nor2_1 _4787_ (.A(net1248),
    .B(_0514_),
    .Y(_0516_));
 sg13g2_xnor2_1 _4788_ (.Y(_0517_),
    .A(net1214),
    .B(_0511_));
 sg13g2_o21ai_1 _4789_ (.B1(_0515_),
    .Y(_0518_),
    .A1(net1262),
    .A2(_0493_));
 sg13g2_nor4_1 _4790_ (.A(_0508_),
    .B(_0516_),
    .C(_0517_),
    .D(_0518_),
    .Y(_0519_));
 sg13g2_or3_1 _4791_ (.A(net1215),
    .B(_0511_),
    .C(_0516_),
    .X(_0520_));
 sg13g2_nand2_1 _4792_ (.Y(_0521_),
    .A(_0515_),
    .B(_0520_));
 sg13g2_nand2b_1 _4793_ (.Y(_0522_),
    .B(_0505_),
    .A_N(_0504_));
 sg13g2_a221oi_1 _4794_ (.B2(_0507_),
    .C1(_0419_),
    .B1(_0521_),
    .A1(_0495_),
    .Y(_0523_),
    .A2(_0519_));
 sg13g2_or2_1 _4795_ (.X(_0524_),
    .B(net1208),
    .A(net308));
 sg13g2_a21oi_1 _4796_ (.A1(_0522_),
    .A2(_0523_),
    .Y(_0059_),
    .B1(_0524_));
 sg13g2_and2_1 _4797_ (.A(net1319),
    .B(net310),
    .X(_0060_));
 sg13g2_o21ai_1 _4798_ (.B1(net1148),
    .Y(_0525_),
    .A1(net1228),
    .A2(net1137));
 sg13g2_nor2b_1 _4799_ (.A(net1228),
    .B_N(net1143),
    .Y(_0526_));
 sg13g2_nor2_2 _4800_ (.A(_0525_),
    .B(_0526_),
    .Y(_0527_));
 sg13g2_a21oi_1 _4801_ (.A1(net1222),
    .A2(net1153),
    .Y(_0528_),
    .B1(net1148));
 sg13g2_nor2_1 _4802_ (.A(_0527_),
    .B(_0528_),
    .Y(_0529_));
 sg13g2_o21ai_1 _4803_ (.B1(_0527_),
    .Y(_0530_),
    .A1(\s0.was_valid_out[15] [0]),
    .A2(net1141));
 sg13g2_nor2_1 _4804_ (.A(net1136),
    .B(_0525_),
    .Y(_0531_));
 sg13g2_o21ai_1 _4805_ (.B1(net923),
    .Y(_0532_),
    .A1(\s0.was_valid_out[15] [0]),
    .A2(net1153));
 sg13g2_nand2_1 _4806_ (.Y(_0533_),
    .A(_0530_),
    .B(_0532_));
 sg13g2_o21ai_1 _4807_ (.B1(net1319),
    .Y(_0534_),
    .A1(_0531_),
    .A2(_0533_));
 sg13g2_a21oi_1 _4808_ (.A1(_2446_),
    .A2(_0529_),
    .Y(_0061_),
    .B1(_0534_));
 sg13g2_nor3_1 _4809_ (.A(net1220),
    .B(_0527_),
    .C(_0528_),
    .Y(_0062_));
 sg13g2_mux2_1 _4810_ (.A0(\s0.data_out[15][0] ),
    .A1(\s0.data_out[16][0] ),
    .S(net1152),
    .X(_0535_));
 sg13g2_nand2_1 _4811_ (.Y(_0536_),
    .A(net922),
    .B(_0535_));
 sg13g2_and2_1 _4812_ (.A(net1134),
    .B(\s0.data_out[15][0] ),
    .X(_0537_));
 sg13g2_nor2b_1 _4813_ (.A(net1134),
    .B_N(net1074),
    .Y(_0538_));
 sg13g2_o21ai_1 _4814_ (.B1(net1149),
    .Y(_0539_),
    .A1(_0537_),
    .A2(_0538_));
 sg13g2_nand3_1 _4815_ (.B(_0536_),
    .C(_0539_),
    .A(net1317),
    .Y(_0540_));
 sg13g2_o21ai_1 _4816_ (.B1(_0540_),
    .Y(_0541_),
    .A1(net1305),
    .A2(net450));
 sg13g2_inv_1 _4817_ (.Y(_0063_),
    .A(_0541_));
 sg13g2_mux2_1 _4818_ (.A0(\s0.data_out[15][1] ),
    .A1(\s0.data_out[16][1] ),
    .S(net1152),
    .X(_0542_));
 sg13g2_nand2_1 _4819_ (.Y(_0543_),
    .A(net922),
    .B(_0542_));
 sg13g2_and2_1 _4820_ (.A(net1135),
    .B(\s0.data_out[15][1] ),
    .X(_0544_));
 sg13g2_nor2b_1 _4821_ (.A(net1135),
    .B_N(net1070),
    .Y(_0545_));
 sg13g2_o21ai_1 _4822_ (.B1(net1149),
    .Y(_0546_),
    .A1(_0544_),
    .A2(_0545_));
 sg13g2_nand3_1 _4823_ (.B(_0543_),
    .C(_0546_),
    .A(net1317),
    .Y(_0547_));
 sg13g2_o21ai_1 _4824_ (.B1(_0547_),
    .Y(_0548_),
    .A1(net1317),
    .A2(net476));
 sg13g2_inv_1 _4825_ (.Y(_0064_),
    .A(_0548_));
 sg13g2_mux2_1 _4826_ (.A0(\s0.data_out[15][2] ),
    .A1(\s0.data_out[16][2] ),
    .S(net1152),
    .X(_0549_));
 sg13g2_nand2_1 _4827_ (.Y(_0550_),
    .A(net922),
    .B(_0549_));
 sg13g2_and2_1 _4828_ (.A(net1134),
    .B(\s0.data_out[15][2] ),
    .X(_0551_));
 sg13g2_nor2b_1 _4829_ (.A(net1134),
    .B_N(net1066),
    .Y(_0552_));
 sg13g2_o21ai_1 _4830_ (.B1(net1149),
    .Y(_0553_),
    .A1(_0551_),
    .A2(_0552_));
 sg13g2_nand3_1 _4831_ (.B(_0550_),
    .C(_0553_),
    .A(net1317),
    .Y(_0554_));
 sg13g2_o21ai_1 _4832_ (.B1(_0554_),
    .Y(_0555_),
    .A1(net1317),
    .A2(net422));
 sg13g2_inv_1 _4833_ (.Y(_0065_),
    .A(_0555_));
 sg13g2_nand2b_1 _4834_ (.Y(_0556_),
    .B(net387),
    .A_N(net1152));
 sg13g2_a21oi_1 _4835_ (.A1(_0489_),
    .A2(_0556_),
    .Y(_0557_),
    .B1(net1149));
 sg13g2_nor2b_1 _4836_ (.A(net1134),
    .B_N(net1062),
    .Y(_0558_));
 sg13g2_a21oi_1 _4837_ (.A1(net1134),
    .A2(net387),
    .Y(_0559_),
    .B1(_0558_));
 sg13g2_o21ai_1 _4838_ (.B1(net1317),
    .Y(_0560_),
    .A1(net922),
    .A2(_0559_));
 sg13g2_nand2_1 _4839_ (.Y(_0561_),
    .A(net1220),
    .B(_2485_));
 sg13g2_o21ai_1 _4840_ (.B1(_0561_),
    .Y(_0562_),
    .A1(_0557_),
    .A2(_0560_));
 sg13g2_inv_1 _4841_ (.Y(_0066_),
    .A(_0562_));
 sg13g2_mux2_1 _4842_ (.A0(\s0.data_out[15][4] ),
    .A1(\s0.data_out[16][4] ),
    .S(net1153),
    .X(_0563_));
 sg13g2_nand2_1 _4843_ (.Y(_0564_),
    .A(net923),
    .B(_0563_));
 sg13g2_and2_1 _4844_ (.A(net1137),
    .B(\s0.data_out[15][4] ),
    .X(_0565_));
 sg13g2_nor2b_1 _4845_ (.A(net1136),
    .B_N(net1059),
    .Y(_0566_));
 sg13g2_o21ai_1 _4846_ (.B1(net1150),
    .Y(_0567_),
    .A1(_0565_),
    .A2(_0566_));
 sg13g2_nand3_1 _4847_ (.B(_0564_),
    .C(_0567_),
    .A(net1319),
    .Y(_0568_));
 sg13g2_o21ai_1 _4848_ (.B1(_0568_),
    .Y(_0569_),
    .A1(net1306),
    .A2(net416));
 sg13g2_inv_1 _4849_ (.Y(_0067_),
    .A(_0569_));
 sg13g2_mux2_1 _4850_ (.A0(\s0.data_out[15][5] ),
    .A1(\s0.data_out[16][5] ),
    .S(net1153),
    .X(_0570_));
 sg13g2_nand2_1 _4851_ (.Y(_0571_),
    .A(net923),
    .B(_0570_));
 sg13g2_and2_1 _4852_ (.A(net1137),
    .B(\s0.data_out[15][5] ),
    .X(_0572_));
 sg13g2_nor2b_1 _4853_ (.A(net1136),
    .B_N(net1055),
    .Y(_0573_));
 sg13g2_o21ai_1 _4854_ (.B1(net1149),
    .Y(_0574_),
    .A1(_0572_),
    .A2(_0573_));
 sg13g2_nand3_1 _4855_ (.B(_0571_),
    .C(_0574_),
    .A(net1323),
    .Y(_0575_));
 sg13g2_o21ai_1 _4856_ (.B1(_0575_),
    .Y(_0576_),
    .A1(net1323),
    .A2(net456));
 sg13g2_inv_1 _4857_ (.Y(_0068_),
    .A(_0576_));
 sg13g2_nand2b_1 _4858_ (.Y(_0577_),
    .B(\s0.data_out[15][6] ),
    .A_N(net1153));
 sg13g2_a21oi_1 _4859_ (.A1(_0496_),
    .A2(_0577_),
    .Y(_0578_),
    .B1(net1148));
 sg13g2_nor2b_1 _4860_ (.A(net1136),
    .B_N(net1051),
    .Y(_0579_));
 sg13g2_a21oi_1 _4861_ (.A1(net1136),
    .A2(\s0.data_out[15][6] ),
    .Y(_0580_),
    .B1(_0579_));
 sg13g2_o21ai_1 _4862_ (.B1(net1317),
    .Y(_0581_),
    .A1(net923),
    .A2(_0580_));
 sg13g2_or2_1 _4863_ (.X(_0582_),
    .B(net546),
    .A(net1318));
 sg13g2_o21ai_1 _4864_ (.B1(_0582_),
    .Y(_0583_),
    .A1(_0578_),
    .A2(_0581_));
 sg13g2_inv_1 _4865_ (.Y(_0069_),
    .A(net547));
 sg13g2_nand2b_1 _4866_ (.Y(_0584_),
    .B(net554),
    .A_N(net1152));
 sg13g2_a21oi_1 _4867_ (.A1(_0500_),
    .A2(_0584_),
    .Y(_0585_),
    .B1(net1149));
 sg13g2_nor2b_1 _4868_ (.A(net1135),
    .B_N(net1047),
    .Y(_0586_));
 sg13g2_a21oi_1 _4869_ (.A1(net1135),
    .A2(net554),
    .Y(_0587_),
    .B1(_0586_));
 sg13g2_o21ai_1 _4870_ (.B1(net1317),
    .Y(_0588_),
    .A1(net922),
    .A2(_0587_));
 sg13g2_or2_1 _4871_ (.X(_0589_),
    .B(net591),
    .A(net1318));
 sg13g2_o21ai_1 _4872_ (.B1(_0589_),
    .Y(_0590_),
    .A1(_0585_),
    .A2(_0588_));
 sg13g2_inv_1 _4873_ (.Y(_0070_),
    .A(_0590_));
 sg13g2_mux2_1 _4874_ (.A0(\s0.data_out[16][2] ),
    .A1(\s0.data_out[15][2] ),
    .S(net1141),
    .X(_0591_));
 sg13g2_a21oi_1 _4875_ (.A1(net1134),
    .A2(_0591_),
    .Y(_0592_),
    .B1(_0552_));
 sg13g2_o21ai_1 _4876_ (.B1(_0550_),
    .Y(_0593_),
    .A1(net922),
    .A2(_0592_));
 sg13g2_mux2_1 _4877_ (.A0(\s0.data_out[16][1] ),
    .A1(\s0.data_out[15][1] ),
    .S(net1141),
    .X(_0594_));
 sg13g2_a21oi_1 _4878_ (.A1(net1135),
    .A2(_0594_),
    .Y(_0595_),
    .B1(_0545_));
 sg13g2_nand2b_1 _4879_ (.Y(_0596_),
    .B(net1149),
    .A_N(_0595_));
 sg13g2_nand3_1 _4880_ (.B(_0543_),
    .C(_0596_),
    .A(net1277),
    .Y(_0597_));
 sg13g2_a21oi_1 _4881_ (.A1(_0543_),
    .A2(_0596_),
    .Y(_0598_),
    .B1(net1277));
 sg13g2_mux2_1 _4882_ (.A0(\s0.data_out[16][0] ),
    .A1(\s0.data_out[15][0] ),
    .S(net1141),
    .X(_0599_));
 sg13g2_a21oi_1 _4883_ (.A1(net1134),
    .A2(_0599_),
    .Y(_0600_),
    .B1(_0538_));
 sg13g2_o21ai_1 _4884_ (.B1(_0536_),
    .Y(_0601_),
    .A1(net922),
    .A2(_0600_));
 sg13g2_nor2b_1 _4885_ (.A(net1282),
    .B_N(_0601_),
    .Y(_0602_));
 sg13g2_a221oi_1 _4886_ (.B2(_0602_),
    .C1(_0598_),
    .B1(_0597_),
    .A1(net1213),
    .Y(_0603_),
    .A2(_0593_));
 sg13g2_nand2_1 _4887_ (.Y(_0604_),
    .A(net1141),
    .B(net387));
 sg13g2_o21ai_1 _4888_ (.B1(_0604_),
    .Y(_0605_),
    .A1(net1141),
    .A2(_2485_));
 sg13g2_a21o_1 _4889_ (.A2(_0605_),
    .A1(net1135),
    .B1(_0558_),
    .X(_0606_));
 sg13g2_a21oi_1 _4890_ (.A1(net1149),
    .A2(_0606_),
    .Y(_0607_),
    .B1(_0557_));
 sg13g2_nand2_1 _4891_ (.Y(_0608_),
    .A(net1264),
    .B(_0607_));
 sg13g2_o21ai_1 _4892_ (.B1(_0608_),
    .Y(_0609_),
    .A1(net1213),
    .A2(_0593_));
 sg13g2_nand2_1 _4893_ (.Y(_0610_),
    .A(net1142),
    .B(net554));
 sg13g2_mux2_1 _4894_ (.A0(\s0.data_out[16][7] ),
    .A1(\s0.data_out[15][7] ),
    .S(net1141),
    .X(_0611_));
 sg13g2_a21o_1 _4895_ (.A2(_0611_),
    .A1(net1136),
    .B1(_0586_),
    .X(_0612_));
 sg13g2_a21oi_1 _4896_ (.A1(net1148),
    .A2(_0612_),
    .Y(_0613_),
    .B1(_0585_));
 sg13g2_nand2_1 _4897_ (.Y(_0614_),
    .A(net1142),
    .B(net562));
 sg13g2_mux2_1 _4898_ (.A0(\s0.data_out[16][6] ),
    .A1(\s0.data_out[15][6] ),
    .S(net1143),
    .X(_0615_));
 sg13g2_a21o_1 _4899_ (.A2(_0615_),
    .A1(net1136),
    .B1(_0579_),
    .X(_0616_));
 sg13g2_a21oi_1 _4900_ (.A1(net1148),
    .A2(_0616_),
    .Y(_0617_),
    .B1(_0578_));
 sg13g2_a22oi_1 _4901_ (.Y(_0618_),
    .B1(_0617_),
    .B2(net1244),
    .A2(_0613_),
    .A1(net1235));
 sg13g2_nor2_1 _4902_ (.A(net1244),
    .B(_0617_),
    .Y(_0619_));
 sg13g2_or2_1 _4903_ (.X(_0620_),
    .B(_0613_),
    .A(net1235));
 sg13g2_nand3b_1 _4904_ (.B(_0620_),
    .C(_0618_),
    .Y(_0621_),
    .A_N(_0619_));
 sg13g2_mux2_1 _4905_ (.A0(\s0.data_out[16][5] ),
    .A1(\s0.data_out[15][5] ),
    .S(net1143),
    .X(_0622_));
 sg13g2_a21oi_1 _4906_ (.A1(net1137),
    .A2(_0622_),
    .Y(_0623_),
    .B1(_0573_));
 sg13g2_nand2b_1 _4907_ (.Y(_0624_),
    .B(net1148),
    .A_N(_0623_));
 sg13g2_a21oi_1 _4908_ (.A1(_0571_),
    .A2(_0624_),
    .Y(_0625_),
    .B1(net1250));
 sg13g2_nand3_1 _4909_ (.B(_0571_),
    .C(_0624_),
    .A(net1250),
    .Y(_0626_));
 sg13g2_mux2_1 _4910_ (.A0(\s0.data_out[16][4] ),
    .A1(\s0.data_out[15][4] ),
    .S(net1141),
    .X(_0627_));
 sg13g2_a21oi_1 _4911_ (.A1(net1136),
    .A2(_0627_),
    .Y(_0628_),
    .B1(_0566_));
 sg13g2_nand2b_1 _4912_ (.Y(_0629_),
    .B(net1148),
    .A_N(_0628_));
 sg13g2_a21oi_1 _4913_ (.A1(_0564_),
    .A2(_0629_),
    .Y(_0630_),
    .B1(net1258));
 sg13g2_nand3_1 _4914_ (.B(_0564_),
    .C(_0629_),
    .A(net1258),
    .Y(_0631_));
 sg13g2_o21ai_1 _4915_ (.B1(_0626_),
    .Y(_0632_),
    .A1(net1264),
    .A2(_0607_));
 sg13g2_nand2b_1 _4916_ (.Y(_0633_),
    .B(_0631_),
    .A_N(_0625_));
 sg13g2_nor4_1 _4917_ (.A(_0621_),
    .B(_0630_),
    .C(_0632_),
    .D(_0633_),
    .Y(_0634_));
 sg13g2_o21ai_1 _4918_ (.B1(_0634_),
    .Y(_0635_),
    .A1(_0603_),
    .A2(_0609_));
 sg13g2_o21ai_1 _4919_ (.B1(_0626_),
    .Y(_0636_),
    .A1(_0625_),
    .A2(_0631_));
 sg13g2_nor2b_1 _4920_ (.A(_0621_),
    .B_N(_0636_),
    .Y(_0637_));
 sg13g2_nor2b_1 _4921_ (.A(_0618_),
    .B_N(_0620_),
    .Y(_0638_));
 sg13g2_nor4_1 _4922_ (.A(_0527_),
    .B(_0528_),
    .C(_0637_),
    .D(_0638_),
    .Y(_0639_));
 sg13g2_or2_1 _4923_ (.X(_0640_),
    .B(net1209),
    .A(net310));
 sg13g2_a21oi_1 _4924_ (.A1(_0635_),
    .A2(_0639_),
    .Y(_0071_),
    .B1(_0640_));
 sg13g2_and2_1 _4925_ (.A(net1319),
    .B(net299),
    .X(_0072_));
 sg13g2_o21ai_1 _4926_ (.B1(net1139),
    .Y(_0641_),
    .A1(net1228),
    .A2(net1125));
 sg13g2_nor2b_1 _4927_ (.A(net1228),
    .B_N(net1130),
    .Y(_0642_));
 sg13g2_nor2_1 _4928_ (.A(_0641_),
    .B(_0642_),
    .Y(_0643_));
 sg13g2_nor2_1 _4929_ (.A(net1140),
    .B(_0526_),
    .Y(_0644_));
 sg13g2_or2_1 _4930_ (.X(_0645_),
    .B(_0644_),
    .A(_0643_));
 sg13g2_or2_1 _4931_ (.X(_0646_),
    .B(net1130),
    .A(net378));
 sg13g2_o21ai_1 _4932_ (.B1(net921),
    .Y(_0647_),
    .A1(net378),
    .A2(net1143));
 sg13g2_o21ai_1 _4933_ (.B1(_0647_),
    .Y(_0648_),
    .A1(net1125),
    .A2(_0641_));
 sg13g2_a21oi_1 _4934_ (.A1(_0643_),
    .A2(_0646_),
    .Y(_0649_),
    .B1(_0648_));
 sg13g2_o21ai_1 _4935_ (.B1(net1319),
    .Y(_0650_),
    .A1(net381),
    .A2(_0645_));
 sg13g2_nor2_1 _4936_ (.A(_0649_),
    .B(_0650_),
    .Y(_0073_));
 sg13g2_nor2_1 _4937_ (.A(net1220),
    .B(_0645_),
    .Y(_0074_));
 sg13g2_mux2_1 _4938_ (.A0(\s0.data_out[14][0] ),
    .A1(\s0.data_out[15][0] ),
    .S(net1142),
    .X(_0651_));
 sg13g2_nand2_1 _4939_ (.Y(_0652_),
    .A(net921),
    .B(_0651_));
 sg13g2_and2_1 _4940_ (.A(net1122),
    .B(\s0.data_out[14][0] ),
    .X(_0653_));
 sg13g2_nor2b_1 _4941_ (.A(net1122),
    .B_N(net1074),
    .Y(_0654_));
 sg13g2_o21ai_1 _4942_ (.B1(net1138),
    .Y(_0655_),
    .A1(_0653_),
    .A2(_0654_));
 sg13g2_nand3_1 _4943_ (.B(_0652_),
    .C(_0655_),
    .A(net1318),
    .Y(_0656_));
 sg13g2_o21ai_1 _4944_ (.B1(_0656_),
    .Y(_0657_),
    .A1(net1318),
    .A2(net461));
 sg13g2_inv_1 _4945_ (.Y(_0075_),
    .A(_0657_));
 sg13g2_mux2_1 _4946_ (.A0(\s0.data_out[14][1] ),
    .A1(\s0.data_out[15][1] ),
    .S(net1142),
    .X(_0658_));
 sg13g2_nand2_1 _4947_ (.Y(_0659_),
    .A(net921),
    .B(_0658_));
 sg13g2_and2_1 _4948_ (.A(net1122),
    .B(\s0.data_out[14][1] ),
    .X(_0660_));
 sg13g2_nor2b_1 _4949_ (.A(net1122),
    .B_N(net1070),
    .Y(_0661_));
 sg13g2_o21ai_1 _4950_ (.B1(net1138),
    .Y(_0662_),
    .A1(_0660_),
    .A2(_0661_));
 sg13g2_nand3_1 _4951_ (.B(_0659_),
    .C(_0662_),
    .A(net1318),
    .Y(_0663_));
 sg13g2_o21ai_1 _4952_ (.B1(_0663_),
    .Y(_0664_),
    .A1(net1318),
    .A2(net431));
 sg13g2_inv_1 _4953_ (.Y(_0076_),
    .A(_0664_));
 sg13g2_mux2_1 _4954_ (.A0(\s0.data_out[14][2] ),
    .A1(\s0.data_out[15][2] ),
    .S(net1142),
    .X(_0665_));
 sg13g2_nand2_1 _4955_ (.Y(_0666_),
    .A(net921),
    .B(_0665_));
 sg13g2_and2_1 _4956_ (.A(net1122),
    .B(\s0.data_out[14][2] ),
    .X(_0667_));
 sg13g2_nor2b_1 _4957_ (.A(net1122),
    .B_N(net1066),
    .Y(_0668_));
 sg13g2_o21ai_1 _4958_ (.B1(net1138),
    .Y(_0669_),
    .A1(_0667_),
    .A2(_0668_));
 sg13g2_nand3_1 _4959_ (.B(_0666_),
    .C(_0669_),
    .A(net1320),
    .Y(_0670_));
 sg13g2_o21ai_1 _4960_ (.B1(_0670_),
    .Y(_0671_),
    .A1(net1320),
    .A2(net445));
 sg13g2_inv_1 _4961_ (.Y(_0077_),
    .A(_0671_));
 sg13g2_o21ai_1 _4962_ (.B1(_0604_),
    .Y(_0672_),
    .A1(net1142),
    .A2(_2486_));
 sg13g2_nand2_1 _4963_ (.Y(_0673_),
    .A(net921),
    .B(_0672_));
 sg13g2_nor2b_1 _4964_ (.A(net1124),
    .B_N(net1063),
    .Y(_0674_));
 sg13g2_a21oi_1 _4965_ (.A1(net1124),
    .A2(net386),
    .Y(_0675_),
    .B1(_0674_));
 sg13g2_o21ai_1 _4966_ (.B1(net1320),
    .Y(_0676_),
    .A1(net921),
    .A2(_0675_));
 sg13g2_nand2b_1 _4967_ (.Y(_0677_),
    .B(_0673_),
    .A_N(_0676_));
 sg13g2_o21ai_1 _4968_ (.B1(_0677_),
    .Y(_0678_),
    .A1(net1320),
    .A2(net387));
 sg13g2_inv_1 _4969_ (.Y(_0078_),
    .A(_0678_));
 sg13g2_mux2_1 _4970_ (.A0(\s0.data_out[14][4] ),
    .A1(\s0.data_out[15][4] ),
    .S(net1143),
    .X(_0679_));
 sg13g2_nand2_1 _4971_ (.Y(_0680_),
    .A(_2464_),
    .B(_0679_));
 sg13g2_and2_1 _4972_ (.A(net1126),
    .B(\s0.data_out[14][4] ),
    .X(_0681_));
 sg13g2_nor2b_1 _4973_ (.A(net1126),
    .B_N(net1059),
    .Y(_0682_));
 sg13g2_o21ai_1 _4974_ (.B1(net1139),
    .Y(_0683_),
    .A1(_0681_),
    .A2(_0682_));
 sg13g2_nand3_1 _4975_ (.B(_0680_),
    .C(_0683_),
    .A(net1322),
    .Y(_0684_));
 sg13g2_o21ai_1 _4976_ (.B1(_0684_),
    .Y(_0685_),
    .A1(net1322),
    .A2(net474));
 sg13g2_inv_1 _4977_ (.Y(_0079_),
    .A(_0685_));
 sg13g2_mux2_1 _4978_ (.A0(\s0.data_out[14][5] ),
    .A1(\s0.data_out[15][5] ),
    .S(net1143),
    .X(_0686_));
 sg13g2_nand2_1 _4979_ (.Y(_0687_),
    .A(_2464_),
    .B(_0686_));
 sg13g2_and2_1 _4980_ (.A(net1125),
    .B(\s0.data_out[14][5] ),
    .X(_0688_));
 sg13g2_nor2b_1 _4981_ (.A(net1125),
    .B_N(net1055),
    .Y(_0689_));
 sg13g2_o21ai_1 _4982_ (.B1(net1139),
    .Y(_0690_),
    .A1(_0688_),
    .A2(_0689_));
 sg13g2_nand3_1 _4983_ (.B(_0687_),
    .C(_0690_),
    .A(net1323),
    .Y(_0691_));
 sg13g2_o21ai_1 _4984_ (.B1(_0691_),
    .Y(_0692_),
    .A1(net1319),
    .A2(net438));
 sg13g2_inv_1 _4985_ (.Y(_0080_),
    .A(_0692_));
 sg13g2_nand2b_1 _4986_ (.Y(_0693_),
    .B(\s0.data_out[14][6] ),
    .A_N(net1142));
 sg13g2_a21oi_1 _4987_ (.A1(_0614_),
    .A2(_0693_),
    .Y(_0694_),
    .B1(net1140));
 sg13g2_nor2b_1 _4988_ (.A(net1125),
    .B_N(net1051),
    .Y(_0695_));
 sg13g2_a21oi_1 _4989_ (.A1(net1125),
    .A2(\s0.data_out[14][6] ),
    .Y(_0696_),
    .B1(_0695_));
 sg13g2_o21ai_1 _4990_ (.B1(net1320),
    .Y(_0697_),
    .A1(net921),
    .A2(_0696_));
 sg13g2_or2_1 _4991_ (.X(_0698_),
    .B(net562),
    .A(net1319));
 sg13g2_o21ai_1 _4992_ (.B1(_0698_),
    .Y(_0699_),
    .A1(_0694_),
    .A2(_0697_));
 sg13g2_inv_1 _4993_ (.Y(_0081_),
    .A(net563));
 sg13g2_nand2b_1 _4994_ (.Y(_0700_),
    .B(\s0.data_out[14][7] ),
    .A_N(net1142));
 sg13g2_a21oi_1 _4995_ (.A1(_0610_),
    .A2(_0700_),
    .Y(_0701_),
    .B1(net1139));
 sg13g2_nor2b_1 _4996_ (.A(net1123),
    .B_N(net1047),
    .Y(_0702_));
 sg13g2_a21oi_1 _4997_ (.A1(net1123),
    .A2(\s0.data_out[14][7] ),
    .Y(_0703_),
    .B1(_0702_));
 sg13g2_o21ai_1 _4998_ (.B1(net1320),
    .Y(_0704_),
    .A1(net921),
    .A2(_0703_));
 sg13g2_or2_1 _4999_ (.X(_0705_),
    .B(net554),
    .A(net1318));
 sg13g2_o21ai_1 _5000_ (.B1(_0705_),
    .Y(_0706_),
    .A1(_0701_),
    .A2(_0704_));
 sg13g2_inv_1 _5001_ (.Y(_0082_),
    .A(net555));
 sg13g2_nand2_1 _5002_ (.Y(_0707_),
    .A(net1131),
    .B(net573));
 sg13g2_mux2_1 _5003_ (.A0(\s0.data_out[15][2] ),
    .A1(\s0.data_out[14][2] ),
    .S(net1130),
    .X(_0708_));
 sg13g2_a21oi_1 _5004_ (.A1(net1123),
    .A2(_0708_),
    .Y(_0709_),
    .B1(_0668_));
 sg13g2_nand2b_1 _5005_ (.Y(_0710_),
    .B(net1138),
    .A_N(_0709_));
 sg13g2_a21o_1 _5006_ (.A2(_0710_),
    .A1(_0666_),
    .B1(net1271),
    .X(_0711_));
 sg13g2_nand2_1 _5007_ (.Y(_0712_),
    .A(net1131),
    .B(net564));
 sg13g2_mux2_1 _5008_ (.A0(\s0.data_out[15][1] ),
    .A1(\s0.data_out[14][1] ),
    .S(net1130),
    .X(_0713_));
 sg13g2_a21oi_1 _5009_ (.A1(net1122),
    .A2(_0713_),
    .Y(_0714_),
    .B1(_0661_));
 sg13g2_nand2b_1 _5010_ (.Y(_0715_),
    .B(net1138),
    .A_N(_0714_));
 sg13g2_and2_1 _5011_ (.A(_0659_),
    .B(_0715_),
    .X(_0716_));
 sg13g2_mux2_1 _5012_ (.A0(\s0.data_out[15][0] ),
    .A1(\s0.data_out[14][0] ),
    .S(net1130),
    .X(_0717_));
 sg13g2_a21oi_1 _5013_ (.A1(net1122),
    .A2(_0717_),
    .Y(_0718_),
    .B1(_0654_));
 sg13g2_nand2b_1 _5014_ (.Y(_0719_),
    .B(net1138),
    .A_N(_0718_));
 sg13g2_a221oi_1 _5015_ (.B2(_0652_),
    .C1(net1282),
    .B1(_0719_),
    .A1(net1277),
    .Y(_0720_),
    .A2(_0716_));
 sg13g2_o21ai_1 _5016_ (.B1(_0711_),
    .Y(_0721_),
    .A1(net1277),
    .A2(_0716_));
 sg13g2_and3_1 _5017_ (.X(_0722_),
    .A(net1271),
    .B(_0666_),
    .C(_0710_));
 sg13g2_mux2_1 _5018_ (.A0(\s0.data_out[15][3] ),
    .A1(\s0.data_out[14][3] ),
    .S(net1130),
    .X(_0723_));
 sg13g2_a21oi_1 _5019_ (.A1(net1124),
    .A2(_0723_),
    .Y(_0724_),
    .B1(_0674_));
 sg13g2_nand2b_1 _5020_ (.Y(_0725_),
    .B(net1138),
    .A_N(_0724_));
 sg13g2_and2_1 _5021_ (.A(_0673_),
    .B(_0725_),
    .X(_0726_));
 sg13g2_a21oi_1 _5022_ (.A1(net1264),
    .A2(_0726_),
    .Y(_0727_),
    .B1(_0722_));
 sg13g2_o21ai_1 _5023_ (.B1(_0727_),
    .Y(_0728_),
    .A1(_0720_),
    .A2(_0721_));
 sg13g2_nand2_1 _5024_ (.Y(_0729_),
    .A(net1131),
    .B(net577));
 sg13g2_mux2_1 _5025_ (.A0(\s0.data_out[15][7] ),
    .A1(\s0.data_out[14][7] ),
    .S(net1130),
    .X(_0730_));
 sg13g2_a21o_1 _5026_ (.A2(_0730_),
    .A1(net1123),
    .B1(_0702_),
    .X(_0731_));
 sg13g2_a21oi_1 _5027_ (.A1(net1139),
    .A2(_0731_),
    .Y(_0732_),
    .B1(_0701_));
 sg13g2_nand2_1 _5028_ (.Y(_0733_),
    .A(net1132),
    .B(net598));
 sg13g2_mux2_1 _5029_ (.A0(\s0.data_out[15][6] ),
    .A1(\s0.data_out[14][6] ),
    .S(net1130),
    .X(_0734_));
 sg13g2_a21o_1 _5030_ (.A2(_0734_),
    .A1(net1125),
    .B1(_0695_),
    .X(_0735_));
 sg13g2_a21oi_1 _5031_ (.A1(net1139),
    .A2(_0735_),
    .Y(_0736_),
    .B1(_0694_));
 sg13g2_a22oi_1 _5032_ (.Y(_0737_),
    .B1(_0736_),
    .B2(net1244),
    .A2(_0732_),
    .A1(net1235));
 sg13g2_or2_1 _5033_ (.X(_0738_),
    .B(_0732_),
    .A(net1235));
 sg13g2_or2_1 _5034_ (.X(_0739_),
    .B(_0736_),
    .A(net1244));
 sg13g2_nand3_1 _5035_ (.B(_0738_),
    .C(_0739_),
    .A(_0737_),
    .Y(_0740_));
 sg13g2_inv_1 _5036_ (.Y(_0741_),
    .A(_0740_));
 sg13g2_nand2_1 _5037_ (.Y(_0742_),
    .A(net1132),
    .B(net525));
 sg13g2_mux2_1 _5038_ (.A0(\s0.data_out[15][4] ),
    .A1(\s0.data_out[14][4] ),
    .S(net1133),
    .X(_0743_));
 sg13g2_a21oi_1 _5039_ (.A1(net1126),
    .A2(_0743_),
    .Y(_0744_),
    .B1(_0682_));
 sg13g2_o21ai_1 _5040_ (.B1(_0680_),
    .Y(_0745_),
    .A1(_2464_),
    .A2(_0744_));
 sg13g2_or2_1 _5041_ (.X(_0746_),
    .B(_0745_),
    .A(net1215));
 sg13g2_nand2_1 _5042_ (.Y(_0747_),
    .A(net1132),
    .B(net548));
 sg13g2_mux2_1 _5043_ (.A0(\s0.data_out[15][5] ),
    .A1(\s0.data_out[14][5] ),
    .S(net1133),
    .X(_0748_));
 sg13g2_a21oi_1 _5044_ (.A1(net1125),
    .A2(_0748_),
    .Y(_0749_),
    .B1(_0689_));
 sg13g2_nand2b_1 _5045_ (.Y(_0750_),
    .B(net1139),
    .A_N(_0749_));
 sg13g2_nand3_1 _5046_ (.B(_0687_),
    .C(_0750_),
    .A(net1250),
    .Y(_0751_));
 sg13g2_nor2_1 _5047_ (.A(net1264),
    .B(_0726_),
    .Y(_0752_));
 sg13g2_a21oi_1 _5048_ (.A1(_0687_),
    .A2(_0750_),
    .Y(_0753_),
    .B1(net1250));
 sg13g2_xnor2_1 _5049_ (.Y(_0754_),
    .A(net1215),
    .B(_0745_));
 sg13g2_nor3_1 _5050_ (.A(_0752_),
    .B(_0753_),
    .C(_0754_),
    .Y(_0755_));
 sg13g2_nand4_1 _5051_ (.B(_0741_),
    .C(_0751_),
    .A(_0728_),
    .Y(_0756_),
    .D(_0755_));
 sg13g2_o21ai_1 _5052_ (.B1(_0751_),
    .Y(_0757_),
    .A1(_0746_),
    .A2(_0753_));
 sg13g2_nor2b_1 _5053_ (.A(_0740_),
    .B_N(_0757_),
    .Y(_0758_));
 sg13g2_nor2b_1 _5054_ (.A(_0737_),
    .B_N(_0738_),
    .Y(_0759_));
 sg13g2_nor3_1 _5055_ (.A(_0645_),
    .B(_0758_),
    .C(_0759_),
    .Y(_0760_));
 sg13g2_or2_1 _5056_ (.X(_0761_),
    .B(net1209),
    .A(net299));
 sg13g2_a21oi_1 _5057_ (.A1(_0756_),
    .A2(_0760_),
    .Y(_0083_),
    .B1(_0761_));
 sg13g2_and2_1 _5058_ (.A(net1321),
    .B(net303),
    .X(_0084_));
 sg13g2_o21ai_1 _5059_ (.B1(net1129),
    .Y(_0762_),
    .A1(net1228),
    .A2(net1114));
 sg13g2_a21oi_1 _5060_ (.A1(_2449_),
    .A2(net1119),
    .Y(_0763_),
    .B1(_0762_));
 sg13g2_inv_1 _5061_ (.Y(_0764_),
    .A(_0763_));
 sg13g2_o21ai_1 _5062_ (.B1(_0764_),
    .Y(_0765_),
    .A1(net1126),
    .A2(_0642_));
 sg13g2_o21ai_1 _5063_ (.B1(_0763_),
    .Y(_0766_),
    .A1(net346),
    .A2(net1119));
 sg13g2_nor2_1 _5064_ (.A(net1114),
    .B(_0762_),
    .Y(_0767_));
 sg13g2_o21ai_1 _5065_ (.B1(net937),
    .Y(_0768_),
    .A1(net346),
    .A2(net1132));
 sg13g2_nor2b_1 _5066_ (.A(_0767_),
    .B_N(_0768_),
    .Y(_0769_));
 sg13g2_o21ai_1 _5067_ (.B1(net1321),
    .Y(_0770_),
    .A1(net378),
    .A2(_0765_));
 sg13g2_a21oi_1 _5068_ (.A1(_0766_),
    .A2(_0769_),
    .Y(_0085_),
    .B1(_0770_));
 sg13g2_nor2_1 _5069_ (.A(net1220),
    .B(_0765_),
    .Y(_0086_));
 sg13g2_mux2_1 _5070_ (.A0(\s0.data_out[13][0] ),
    .A1(\s0.data_out[14][0] ),
    .S(net1131),
    .X(_0771_));
 sg13g2_nand2_1 _5071_ (.Y(_0772_),
    .A(net937),
    .B(_0771_));
 sg13g2_and2_1 _5072_ (.A(net1113),
    .B(\s0.data_out[13][0] ),
    .X(_0773_));
 sg13g2_nor2b_1 _5073_ (.A(net1113),
    .B_N(net1075),
    .Y(_0774_));
 sg13g2_o21ai_1 _5074_ (.B1(net1127),
    .Y(_0775_),
    .A1(_0773_),
    .A2(_0774_));
 sg13g2_nand3_1 _5075_ (.B(_0772_),
    .C(_0775_),
    .A(net1321),
    .Y(_0776_));
 sg13g2_o21ai_1 _5076_ (.B1(_0776_),
    .Y(_0777_),
    .A1(net1321),
    .A2(net457));
 sg13g2_inv_1 _5077_ (.Y(_0087_),
    .A(_0777_));
 sg13g2_nand2b_1 _5078_ (.Y(_0778_),
    .B(net471),
    .A_N(net1131));
 sg13g2_a21oi_1 _5079_ (.A1(_0712_),
    .A2(_0778_),
    .Y(_0779_),
    .B1(net1127));
 sg13g2_nor2b_1 _5080_ (.A(net1112),
    .B_N(net1070),
    .Y(_0780_));
 sg13g2_a21oi_1 _5081_ (.A1(net1112),
    .A2(net471),
    .Y(_0781_),
    .B1(_0780_));
 sg13g2_o21ai_1 _5082_ (.B1(net1333),
    .Y(_0782_),
    .A1(net937),
    .A2(_0781_));
 sg13g2_or2_1 _5083_ (.X(_0783_),
    .B(net564),
    .A(net1320));
 sg13g2_o21ai_1 _5084_ (.B1(_0783_),
    .Y(_0784_),
    .A1(_0779_),
    .A2(_0782_));
 sg13g2_inv_1 _5085_ (.Y(_0088_),
    .A(_0784_));
 sg13g2_nand2b_1 _5086_ (.Y(_0785_),
    .B(net477),
    .A_N(net1131));
 sg13g2_a21oi_1 _5087_ (.A1(_0707_),
    .A2(_0785_),
    .Y(_0786_),
    .B1(net1127));
 sg13g2_nor2b_1 _5088_ (.A(net1112),
    .B_N(net1066),
    .Y(_0787_));
 sg13g2_a21oi_1 _5089_ (.A1(net1112),
    .A2(net477),
    .Y(_0788_),
    .B1(_0787_));
 sg13g2_o21ai_1 _5090_ (.B1(net1333),
    .Y(_0789_),
    .A1(net937),
    .A2(_0788_));
 sg13g2_or2_1 _5091_ (.X(_0790_),
    .B(net573),
    .A(net1333));
 sg13g2_o21ai_1 _5092_ (.B1(_0790_),
    .Y(_0791_),
    .A1(_0786_),
    .A2(_0789_));
 sg13g2_inv_1 _5093_ (.Y(_0089_),
    .A(_0791_));
 sg13g2_mux2_1 _5094_ (.A0(\s0.data_out[13][3] ),
    .A1(\s0.data_out[14][3] ),
    .S(net1131),
    .X(_0792_));
 sg13g2_nand2_1 _5095_ (.Y(_0793_),
    .A(net937),
    .B(_0792_));
 sg13g2_and2_1 _5096_ (.A(net1113),
    .B(\s0.data_out[13][3] ),
    .X(_0794_));
 sg13g2_nor2b_1 _5097_ (.A(net1113),
    .B_N(net1063),
    .Y(_0795_));
 sg13g2_o21ai_1 _5098_ (.B1(net1127),
    .Y(_0796_),
    .A1(_0794_),
    .A2(_0795_));
 sg13g2_nand3_1 _5099_ (.B(_0793_),
    .C(_0796_),
    .A(net1321),
    .Y(_0797_));
 sg13g2_o21ai_1 _5100_ (.B1(_0797_),
    .Y(_0798_),
    .A1(net1320),
    .A2(net386));
 sg13g2_inv_1 _5101_ (.Y(_0090_),
    .A(_0798_));
 sg13g2_nand2b_1 _5102_ (.Y(_0799_),
    .B(net430),
    .A_N(net1132));
 sg13g2_a21oi_1 _5103_ (.A1(_0742_),
    .A2(_0799_),
    .Y(_0800_),
    .B1(net1128));
 sg13g2_nor2b_1 _5104_ (.A(net1115),
    .B_N(net1060),
    .Y(_0801_));
 sg13g2_a21oi_1 _5105_ (.A1(net1115),
    .A2(net430),
    .Y(_0802_),
    .B1(_0801_));
 sg13g2_o21ai_1 _5106_ (.B1(net1322),
    .Y(_0803_),
    .A1(_2452_),
    .A2(_0802_));
 sg13g2_or2_1 _5107_ (.X(_0804_),
    .B(net525),
    .A(net1322));
 sg13g2_o21ai_1 _5108_ (.B1(_0804_),
    .Y(_0805_),
    .A1(_0800_),
    .A2(_0803_));
 sg13g2_inv_1 _5109_ (.Y(_0091_),
    .A(_0805_));
 sg13g2_nand2b_1 _5110_ (.Y(_0806_),
    .B(\s0.data_out[13][5] ),
    .A_N(net1132));
 sg13g2_a21oi_1 _5111_ (.A1(_0747_),
    .A2(_0806_),
    .Y(_0807_),
    .B1(net1128));
 sg13g2_nor2b_1 _5112_ (.A(net1114),
    .B_N(net1056),
    .Y(_0808_));
 sg13g2_a21oi_1 _5113_ (.A1(net1114),
    .A2(\s0.data_out[13][5] ),
    .Y(_0809_),
    .B1(_0808_));
 sg13g2_o21ai_1 _5114_ (.B1(net1322),
    .Y(_0810_),
    .A1(net937),
    .A2(_0809_));
 sg13g2_or2_1 _5115_ (.X(_0811_),
    .B(net548),
    .A(net1322));
 sg13g2_o21ai_1 _5116_ (.B1(_0811_),
    .Y(_0812_),
    .A1(_0807_),
    .A2(_0810_));
 sg13g2_inv_1 _5117_ (.Y(_0092_),
    .A(net549));
 sg13g2_nand2b_1 _5118_ (.Y(_0813_),
    .B(net597),
    .A_N(net1132));
 sg13g2_a21oi_1 _5119_ (.A1(_0733_),
    .A2(_0813_),
    .Y(_0814_),
    .B1(net1128));
 sg13g2_nor2b_1 _5120_ (.A(net1115),
    .B_N(net1052),
    .Y(_0815_));
 sg13g2_a21oi_1 _5121_ (.A1(net1114),
    .A2(net597),
    .Y(_0816_),
    .B1(_0815_));
 sg13g2_o21ai_1 _5122_ (.B1(net1333),
    .Y(_0817_),
    .A1(net937),
    .A2(_0816_));
 sg13g2_or2_1 _5123_ (.X(_0818_),
    .B(net598),
    .A(net1321));
 sg13g2_o21ai_1 _5124_ (.B1(_0818_),
    .Y(_0819_),
    .A1(_0814_),
    .A2(_0817_));
 sg13g2_inv_1 _5125_ (.Y(_0093_),
    .A(_0819_));
 sg13g2_nand2b_1 _5126_ (.Y(_0820_),
    .B(\s0.data_out[13][7] ),
    .A_N(net1131));
 sg13g2_a21oi_1 _5127_ (.A1(_0729_),
    .A2(_0820_),
    .Y(_0821_),
    .B1(net1128));
 sg13g2_nor2b_1 _5128_ (.A(net1113),
    .B_N(net1048),
    .Y(_0822_));
 sg13g2_a21oi_1 _5129_ (.A1(net1112),
    .A2(\s0.data_out[13][7] ),
    .Y(_0823_),
    .B1(_0822_));
 sg13g2_o21ai_1 _5130_ (.B1(net1333),
    .Y(_0824_),
    .A1(net937),
    .A2(_0823_));
 sg13g2_or2_1 _5131_ (.X(_0825_),
    .B(net577),
    .A(net1333));
 sg13g2_o21ai_1 _5132_ (.B1(_0825_),
    .Y(_0826_),
    .A1(_0821_),
    .A2(_0824_));
 sg13g2_inv_1 _5133_ (.Y(_0094_),
    .A(net578));
 sg13g2_mux2_1 _5134_ (.A0(\s0.data_out[14][2] ),
    .A1(\s0.data_out[13][2] ),
    .S(net1119),
    .X(_0827_));
 sg13g2_a21o_1 _5135_ (.A2(_0827_),
    .A1(net1112),
    .B1(_0787_),
    .X(_0828_));
 sg13g2_a21oi_1 _5136_ (.A1(net1127),
    .A2(_0828_),
    .Y(_0829_),
    .B1(_0786_));
 sg13g2_nor2_1 _5137_ (.A(net1270),
    .B(_0829_),
    .Y(_0830_));
 sg13g2_mux2_1 _5138_ (.A0(\s0.data_out[14][1] ),
    .A1(\s0.data_out[13][1] ),
    .S(net1119),
    .X(_0831_));
 sg13g2_a21o_1 _5139_ (.A2(_0831_),
    .A1(net1112),
    .B1(_0780_),
    .X(_0832_));
 sg13g2_a21oi_1 _5140_ (.A1(net1127),
    .A2(_0832_),
    .Y(_0833_),
    .B1(_0779_));
 sg13g2_mux2_1 _5141_ (.A0(\s0.data_out[14][0] ),
    .A1(\s0.data_out[13][0] ),
    .S(net1119),
    .X(_0834_));
 sg13g2_a21oi_1 _5142_ (.A1(net1113),
    .A2(_0834_),
    .Y(_0835_),
    .B1(_0774_));
 sg13g2_nand2b_1 _5143_ (.Y(_0836_),
    .B(net1127),
    .A_N(_0835_));
 sg13g2_nor2_1 _5144_ (.A(net1279),
    .B(_0833_),
    .Y(_0837_));
 sg13g2_a221oi_1 _5145_ (.B2(_0772_),
    .C1(net1283),
    .B1(_0836_),
    .A1(net1279),
    .Y(_0838_),
    .A2(_0833_));
 sg13g2_nor3_1 _5146_ (.A(_0830_),
    .B(_0837_),
    .C(_0838_),
    .Y(_0839_));
 sg13g2_nand2_1 _5147_ (.Y(_0840_),
    .A(net1120),
    .B(net507));
 sg13g2_o21ai_1 _5148_ (.B1(_0840_),
    .Y(_0841_),
    .A1(net1119),
    .A2(_2486_));
 sg13g2_a21oi_1 _5149_ (.A1(net1113),
    .A2(_0841_),
    .Y(_0842_),
    .B1(_0795_));
 sg13g2_nand2b_1 _5150_ (.Y(_0843_),
    .B(net1127),
    .A_N(_0842_));
 sg13g2_and2_1 _5151_ (.A(_0793_),
    .B(_0843_),
    .X(_0844_));
 sg13g2_a221oi_1 _5152_ (.B2(net1265),
    .C1(_0839_),
    .B1(_0844_),
    .A1(net1270),
    .Y(_0845_),
    .A2(_0829_));
 sg13g2_nand2_1 _5153_ (.Y(_0846_),
    .A(net1121),
    .B(net584));
 sg13g2_mux2_1 _5154_ (.A0(\s0.data_out[14][7] ),
    .A1(\s0.data_out[13][7] ),
    .S(net1119),
    .X(_0847_));
 sg13g2_a21o_1 _5155_ (.A2(_0847_),
    .A1(net1112),
    .B1(_0822_),
    .X(_0848_));
 sg13g2_a21oi_1 _5156_ (.A1(net1128),
    .A2(_0848_),
    .Y(_0849_),
    .B1(_0821_));
 sg13g2_nand2_1 _5157_ (.Y(_0850_),
    .A(net1121),
    .B(net597));
 sg13g2_mux2_1 _5158_ (.A0(\s0.data_out[14][6] ),
    .A1(\s0.data_out[13][6] ),
    .S(net1120),
    .X(_0851_));
 sg13g2_a21o_1 _5159_ (.A2(_0851_),
    .A1(net1114),
    .B1(_0815_),
    .X(_0852_));
 sg13g2_a21oi_1 _5160_ (.A1(net1128),
    .A2(_0852_),
    .Y(_0853_),
    .B1(_0814_));
 sg13g2_a22oi_1 _5161_ (.Y(_0854_),
    .B1(_0853_),
    .B2(net1242),
    .A2(_0849_),
    .A1(net1236));
 sg13g2_or2_1 _5162_ (.X(_0855_),
    .B(_0849_),
    .A(net1236));
 sg13g2_or2_1 _5163_ (.X(_0856_),
    .B(_0853_),
    .A(net1242));
 sg13g2_nand3_1 _5164_ (.B(_0855_),
    .C(_0856_),
    .A(_0854_),
    .Y(_0857_));
 sg13g2_mux2_1 _5165_ (.A0(\s0.data_out[14][4] ),
    .A1(\s0.data_out[13][4] ),
    .S(net1120),
    .X(_0858_));
 sg13g2_a21o_1 _5166_ (.A2(_0858_),
    .A1(net1115),
    .B1(_0801_),
    .X(_0859_));
 sg13g2_a21oi_1 _5167_ (.A1(net1129),
    .A2(_0859_),
    .Y(_0860_),
    .B1(_0800_));
 sg13g2_nand2_1 _5168_ (.Y(_0861_),
    .A(net1256),
    .B(_0860_));
 sg13g2_nand2_1 _5169_ (.Y(_0862_),
    .A(net1121),
    .B(net599));
 sg13g2_mux2_1 _5170_ (.A0(\s0.data_out[14][5] ),
    .A1(\s0.data_out[13][5] ),
    .S(net1120),
    .X(_0863_));
 sg13g2_a21o_1 _5171_ (.A2(_0863_),
    .A1(net1114),
    .B1(_0808_),
    .X(_0864_));
 sg13g2_a21oi_1 _5172_ (.A1(net1129),
    .A2(_0864_),
    .Y(_0865_),
    .B1(_0807_));
 sg13g2_nor2_1 _5173_ (.A(net1251),
    .B(_0865_),
    .Y(_0866_));
 sg13g2_or2_1 _5174_ (.X(_0867_),
    .B(_0865_),
    .A(net1251));
 sg13g2_or2_1 _5175_ (.X(_0868_),
    .B(_0860_),
    .A(net1256));
 sg13g2_o21ai_1 _5176_ (.B1(_0868_),
    .Y(_0869_),
    .A1(net1265),
    .A2(_0844_));
 sg13g2_nand2_1 _5177_ (.Y(_0870_),
    .A(net1251),
    .B(_0865_));
 sg13g2_nand3_1 _5178_ (.B(_0867_),
    .C(_0870_),
    .A(_0861_),
    .Y(_0871_));
 sg13g2_or4_1 _5179_ (.A(_0845_),
    .B(_0857_),
    .C(_0869_),
    .D(_0871_),
    .X(_0872_));
 sg13g2_o21ai_1 _5180_ (.B1(_0870_),
    .Y(_0873_),
    .A1(_0861_),
    .A2(_0866_));
 sg13g2_nor2b_1 _5181_ (.A(_0857_),
    .B_N(_0873_),
    .Y(_0874_));
 sg13g2_nor2b_1 _5182_ (.A(_0854_),
    .B_N(_0855_),
    .Y(_0875_));
 sg13g2_nor3_1 _5183_ (.A(_0765_),
    .B(_0874_),
    .C(_0875_),
    .Y(_0876_));
 sg13g2_or2_1 _5184_ (.X(_0877_),
    .B(net1209),
    .A(net303));
 sg13g2_a21oi_1 _5185_ (.A1(_0872_),
    .A2(_0876_),
    .Y(_0095_),
    .B1(_0877_));
 sg13g2_and2_1 _5186_ (.A(net1338),
    .B(net298),
    .X(_0096_));
 sg13g2_o21ai_1 _5187_ (.B1(net1117),
    .Y(_0878_),
    .A1(net1229),
    .A2(net1106));
 sg13g2_nor2b_1 _5188_ (.A(net1229),
    .B_N(net1110),
    .Y(_0879_));
 sg13g2_nor2_1 _5189_ (.A(_0878_),
    .B(_0879_),
    .Y(_0880_));
 sg13g2_a21oi_1 _5190_ (.A1(_2449_),
    .A2(net1119),
    .Y(_0881_),
    .B1(net1114));
 sg13g2_nor2_1 _5191_ (.A(_0880_),
    .B(_0881_),
    .Y(_0882_));
 sg13g2_o21ai_1 _5192_ (.B1(_0880_),
    .Y(_0883_),
    .A1(\s0.was_valid_out[12] [0]),
    .A2(net1111));
 sg13g2_nor2_1 _5193_ (.A(net1107),
    .B(_0878_),
    .Y(_0884_));
 sg13g2_o21ai_1 _5194_ (.B1(net936),
    .Y(_0885_),
    .A1(\s0.was_valid_out[12] [0]),
    .A2(\s0.valid_out[13] [0]));
 sg13g2_nand2_1 _5195_ (.Y(_0886_),
    .A(_0883_),
    .B(_0885_));
 sg13g2_o21ai_1 _5196_ (.B1(net1338),
    .Y(_0887_),
    .A1(_0884_),
    .A2(_0886_));
 sg13g2_a21oi_1 _5197_ (.A1(_2445_),
    .A2(_0882_),
    .Y(_0097_),
    .B1(_0887_));
 sg13g2_nor3_1 _5198_ (.A(net1220),
    .B(_0880_),
    .C(_0881_),
    .Y(_0098_));
 sg13g2_mux2_1 _5199_ (.A0(\s0.data_out[12][0] ),
    .A1(\s0.data_out[13][0] ),
    .S(net1120),
    .X(_0888_));
 sg13g2_nand2_1 _5200_ (.Y(_0889_),
    .A(net935),
    .B(_0888_));
 sg13g2_and2_1 _5201_ (.A(net1100),
    .B(\s0.data_out[12][0] ),
    .X(_0890_));
 sg13g2_nor2b_1 _5202_ (.A(net1100),
    .B_N(net1075),
    .Y(_0891_));
 sg13g2_o21ai_1 _5203_ (.B1(net1116),
    .Y(_0892_),
    .A1(_0890_),
    .A2(_0891_));
 sg13g2_nand3_1 _5204_ (.B(_0889_),
    .C(_0892_),
    .A(net1332),
    .Y(_0893_));
 sg13g2_o21ai_1 _5205_ (.B1(_0893_),
    .Y(_0894_),
    .A1(net1333),
    .A2(net439));
 sg13g2_inv_1 _5206_ (.Y(_0099_),
    .A(_0894_));
 sg13g2_mux2_1 _5207_ (.A0(\s0.data_out[12][1] ),
    .A1(\s0.data_out[13][1] ),
    .S(net1120),
    .X(_0895_));
 sg13g2_nand2_1 _5208_ (.Y(_0896_),
    .A(net935),
    .B(_0895_));
 sg13g2_and2_1 _5209_ (.A(net1100),
    .B(\s0.data_out[12][1] ),
    .X(_0897_));
 sg13g2_nor2b_1 _5210_ (.A(net1100),
    .B_N(net1070),
    .Y(_0898_));
 sg13g2_o21ai_1 _5211_ (.B1(net1116),
    .Y(_0899_),
    .A1(_0897_),
    .A2(_0898_));
 sg13g2_nand3_1 _5212_ (.B(_0896_),
    .C(_0899_),
    .A(net1332),
    .Y(_0900_));
 sg13g2_o21ai_1 _5213_ (.B1(_0900_),
    .Y(_0901_),
    .A1(net1332),
    .A2(net471));
 sg13g2_inv_1 _5214_ (.Y(_0100_),
    .A(_0901_));
 sg13g2_mux2_1 _5215_ (.A0(\s0.data_out[12][2] ),
    .A1(\s0.data_out[13][2] ),
    .S(net1121),
    .X(_0902_));
 sg13g2_nand2_1 _5216_ (.Y(_0903_),
    .A(net935),
    .B(_0902_));
 sg13g2_and2_1 _5217_ (.A(net1100),
    .B(net612),
    .X(_0904_));
 sg13g2_nor2b_1 _5218_ (.A(net1101),
    .B_N(net1066),
    .Y(_0905_));
 sg13g2_o21ai_1 _5219_ (.B1(net1117),
    .Y(_0906_),
    .A1(_0904_),
    .A2(_0905_));
 sg13g2_nand3_1 _5220_ (.B(_0903_),
    .C(_0906_),
    .A(net1332),
    .Y(_0907_));
 sg13g2_o21ai_1 _5221_ (.B1(_0907_),
    .Y(_0908_),
    .A1(net1332),
    .A2(net477));
 sg13g2_inv_1 _5222_ (.Y(_0101_),
    .A(_0908_));
 sg13g2_nand2b_1 _5223_ (.Y(_0909_),
    .B(net472),
    .A_N(net1121));
 sg13g2_a21oi_1 _5224_ (.A1(_0840_),
    .A2(_0909_),
    .Y(_0910_),
    .B1(net1117));
 sg13g2_nor2b_1 _5225_ (.A(net1101),
    .B_N(net1063),
    .Y(_0911_));
 sg13g2_a21oi_1 _5226_ (.A1(net1101),
    .A2(net472),
    .Y(_0912_),
    .B1(_0911_));
 sg13g2_o21ai_1 _5227_ (.B1(net1332),
    .Y(_0913_),
    .A1(net935),
    .A2(_0912_));
 sg13g2_or2_1 _5228_ (.X(_0914_),
    .B(net507),
    .A(net1332));
 sg13g2_o21ai_1 _5229_ (.B1(_0914_),
    .Y(_0915_),
    .A1(_0910_),
    .A2(_0913_));
 sg13g2_inv_1 _5230_ (.Y(_0102_),
    .A(net508));
 sg13g2_mux2_1 _5231_ (.A0(\s0.data_out[12][4] ),
    .A1(\s0.data_out[13][4] ),
    .S(net1120),
    .X(_0916_));
 sg13g2_nand2_1 _5232_ (.Y(_0917_),
    .A(net935),
    .B(_0916_));
 sg13g2_and2_1 _5233_ (.A(net1102),
    .B(\s0.data_out[12][4] ),
    .X(_0918_));
 sg13g2_nor2b_1 _5234_ (.A(net1102),
    .B_N(net1060),
    .Y(_0919_));
 sg13g2_o21ai_1 _5235_ (.B1(net1116),
    .Y(_0920_),
    .A1(_0918_),
    .A2(_0919_));
 sg13g2_nand3_1 _5236_ (.B(_0917_),
    .C(_0920_),
    .A(net1334),
    .Y(_0921_));
 sg13g2_o21ai_1 _5237_ (.B1(_0921_),
    .Y(_0922_),
    .A1(net1334),
    .A2(net430));
 sg13g2_inv_1 _5238_ (.Y(_0103_),
    .A(_0922_));
 sg13g2_nand2b_1 _5239_ (.Y(_0923_),
    .B(net501),
    .A_N(net1121));
 sg13g2_a21oi_1 _5240_ (.A1(_0862_),
    .A2(_0923_),
    .Y(_0924_),
    .B1(net1117));
 sg13g2_nor2b_1 _5241_ (.A(net1106),
    .B_N(net1056),
    .Y(_0925_));
 sg13g2_a21oi_1 _5242_ (.A1(net1106),
    .A2(net501),
    .Y(_0926_),
    .B1(_0925_));
 sg13g2_o21ai_1 _5243_ (.B1(net1338),
    .Y(_0927_),
    .A1(net936),
    .A2(_0926_));
 sg13g2_or2_1 _5244_ (.X(_0928_),
    .B(net599),
    .A(net1338));
 sg13g2_o21ai_1 _5245_ (.B1(_0928_),
    .Y(_0929_),
    .A1(_0924_),
    .A2(_0927_));
 sg13g2_inv_1 _5246_ (.Y(_0104_),
    .A(_0929_));
 sg13g2_nand2b_1 _5247_ (.Y(_0930_),
    .B(net588),
    .A_N(net1121));
 sg13g2_a21oi_1 _5248_ (.A1(_0850_),
    .A2(_0930_),
    .Y(_0931_),
    .B1(net1117));
 sg13g2_nor2b_1 _5249_ (.A(net1107),
    .B_N(net1052),
    .Y(_0932_));
 sg13g2_a21oi_1 _5250_ (.A1(net1107),
    .A2(net588),
    .Y(_0933_),
    .B1(_0932_));
 sg13g2_o21ai_1 _5251_ (.B1(net1338),
    .Y(_0934_),
    .A1(net936),
    .A2(_0933_));
 sg13g2_or2_1 _5252_ (.X(_0935_),
    .B(net597),
    .A(net1338));
 sg13g2_o21ai_1 _5253_ (.B1(_0935_),
    .Y(_0936_),
    .A1(_0931_),
    .A2(_0934_));
 sg13g2_inv_1 _5254_ (.Y(_0105_),
    .A(_0936_));
 sg13g2_nand2b_1 _5255_ (.Y(_0937_),
    .B(\s0.data_out[12][7] ),
    .A_N(net1121));
 sg13g2_a21oi_1 _5256_ (.A1(_0846_),
    .A2(_0937_),
    .Y(_0938_),
    .B1(net1118));
 sg13g2_nor2b_1 _5257_ (.A(net1107),
    .B_N(net1048),
    .Y(_0939_));
 sg13g2_a21oi_1 _5258_ (.A1(net1107),
    .A2(\s0.data_out[12][7] ),
    .Y(_0940_),
    .B1(_0939_));
 sg13g2_o21ai_1 _5259_ (.B1(net1338),
    .Y(_0941_),
    .A1(net936),
    .A2(_0940_));
 sg13g2_or2_1 _5260_ (.X(_0942_),
    .B(net584),
    .A(net1338));
 sg13g2_o21ai_1 _5261_ (.B1(_0942_),
    .Y(_0943_),
    .A1(_0938_),
    .A2(_0941_));
 sg13g2_inv_1 _5262_ (.Y(_0106_),
    .A(net585));
 sg13g2_nand2_1 _5263_ (.Y(_0944_),
    .A(net1108),
    .B(net504));
 sg13g2_o21ai_1 _5264_ (.B1(_0944_),
    .Y(_0945_),
    .A1(net1108),
    .A2(_2487_));
 sg13g2_a21oi_1 _5265_ (.A1(net1101),
    .A2(_0945_),
    .Y(_0946_),
    .B1(_0905_));
 sg13g2_o21ai_1 _5266_ (.B1(_0903_),
    .Y(_0947_),
    .A1(net935),
    .A2(_0946_));
 sg13g2_nand2_1 _5267_ (.Y(_0948_),
    .A(net1109),
    .B(net528));
 sg13g2_mux2_1 _5268_ (.A0(\s0.data_out[13][1] ),
    .A1(\s0.data_out[12][1] ),
    .S(net1108),
    .X(_0949_));
 sg13g2_a21oi_1 _5269_ (.A1(net1100),
    .A2(_0949_),
    .Y(_0950_),
    .B1(_0898_));
 sg13g2_nand2b_1 _5270_ (.Y(_0951_),
    .B(net1116),
    .A_N(_0950_));
 sg13g2_nand3_1 _5271_ (.B(_0896_),
    .C(_0951_),
    .A(net1279),
    .Y(_0952_));
 sg13g2_mux2_1 _5272_ (.A0(\s0.data_out[13][0] ),
    .A1(\s0.data_out[12][0] ),
    .S(net1108),
    .X(_0953_));
 sg13g2_a21oi_1 _5273_ (.A1(net1100),
    .A2(_0953_),
    .Y(_0954_),
    .B1(_0891_));
 sg13g2_o21ai_1 _5274_ (.B1(_0889_),
    .Y(_0955_),
    .A1(net935),
    .A2(_0954_));
 sg13g2_nor2b_1 _5275_ (.A(net1282),
    .B_N(_0955_),
    .Y(_0956_));
 sg13g2_a21oi_1 _5276_ (.A1(_0896_),
    .A2(_0951_),
    .Y(_0957_),
    .B1(net1279));
 sg13g2_a221oi_1 _5277_ (.B2(_0956_),
    .C1(_0957_),
    .B1(_0952_),
    .A1(net1212),
    .Y(_0958_),
    .A2(_0947_));
 sg13g2_mux2_1 _5278_ (.A0(\s0.data_out[13][3] ),
    .A1(\s0.data_out[12][3] ),
    .S(net1108),
    .X(_0959_));
 sg13g2_a21o_1 _5279_ (.A2(_0959_),
    .A1(net1100),
    .B1(_0911_),
    .X(_0960_));
 sg13g2_a21oi_1 _5280_ (.A1(net1117),
    .A2(_0960_),
    .Y(_0961_),
    .B1(_0910_));
 sg13g2_nand2_1 _5281_ (.Y(_0962_),
    .A(net1265),
    .B(_0961_));
 sg13g2_or2_1 _5282_ (.X(_0963_),
    .B(_0947_),
    .A(net1212));
 sg13g2_nand3b_1 _5283_ (.B(_0962_),
    .C(_0963_),
    .Y(_0964_),
    .A_N(_0958_));
 sg13g2_nand2_1 _5284_ (.Y(_0965_),
    .A(net1110),
    .B(net594));
 sg13g2_mux2_1 _5285_ (.A0(\s0.data_out[13][7] ),
    .A1(\s0.data_out[12][7] ),
    .S(net1111),
    .X(_0966_));
 sg13g2_a21o_1 _5286_ (.A2(_0966_),
    .A1(net1107),
    .B1(_0939_),
    .X(_0967_));
 sg13g2_a21oi_1 _5287_ (.A1(net1117),
    .A2(_0967_),
    .Y(_0968_),
    .B1(_0938_));
 sg13g2_nand2_1 _5288_ (.Y(_0969_),
    .A(net1111),
    .B(net588));
 sg13g2_mux2_1 _5289_ (.A0(\s0.data_out[13][6] ),
    .A1(\s0.data_out[12][6] ),
    .S(net1111),
    .X(_0970_));
 sg13g2_a21o_1 _5290_ (.A2(_0970_),
    .A1(net1107),
    .B1(_0932_),
    .X(_0971_));
 sg13g2_a21oi_1 _5291_ (.A1(net1118),
    .A2(_0971_),
    .Y(_0972_),
    .B1(_0931_));
 sg13g2_a22oi_1 _5292_ (.Y(_0973_),
    .B1(_0972_),
    .B2(net1242),
    .A2(_0968_),
    .A1(net1236));
 sg13g2_or2_1 _5293_ (.X(_0974_),
    .B(_0972_),
    .A(net1242));
 sg13g2_nor2_1 _5294_ (.A(net1236),
    .B(_0968_),
    .Y(_0975_));
 sg13g2_or2_1 _5295_ (.X(_0976_),
    .B(_0968_),
    .A(net1236));
 sg13g2_and3_1 _5296_ (.X(_0977_),
    .A(_0973_),
    .B(_0974_),
    .C(_0976_));
 sg13g2_nand2_1 _5297_ (.Y(_0978_),
    .A(net1109),
    .B(\s0.data_out[12][4] ));
 sg13g2_mux2_1 _5298_ (.A0(\s0.data_out[13][4] ),
    .A1(\s0.data_out[12][4] ),
    .S(net1108),
    .X(_0979_));
 sg13g2_a21oi_1 _5299_ (.A1(net1102),
    .A2(_0979_),
    .Y(_0980_),
    .B1(_0919_));
 sg13g2_o21ai_1 _5300_ (.B1(_0917_),
    .Y(_0981_),
    .A1(net935),
    .A2(_0980_));
 sg13g2_or2_1 _5301_ (.X(_0982_),
    .B(_0981_),
    .A(net1215));
 sg13g2_nand2_1 _5302_ (.Y(_0983_),
    .A(net1111),
    .B(net501));
 sg13g2_mux2_1 _5303_ (.A0(\s0.data_out[13][5] ),
    .A1(\s0.data_out[12][5] ),
    .S(net1110),
    .X(_0984_));
 sg13g2_a21o_1 _5304_ (.A2(_0984_),
    .A1(net1106),
    .B1(_0925_),
    .X(_0985_));
 sg13g2_a21oi_1 _5305_ (.A1(net1117),
    .A2(_0985_),
    .Y(_0986_),
    .B1(_0924_));
 sg13g2_nand2_1 _5306_ (.Y(_0987_),
    .A(net1251),
    .B(_0986_));
 sg13g2_nor2_1 _5307_ (.A(net1251),
    .B(_0986_),
    .Y(_0988_));
 sg13g2_nor2_1 _5308_ (.A(net1265),
    .B(_0961_),
    .Y(_0989_));
 sg13g2_xnor2_1 _5309_ (.Y(_0990_),
    .A(net1215),
    .B(_0981_));
 sg13g2_nor3_1 _5310_ (.A(_0988_),
    .B(_0989_),
    .C(_0990_),
    .Y(_0991_));
 sg13g2_and3_1 _5311_ (.X(_0992_),
    .A(_0977_),
    .B(_0987_),
    .C(_0991_));
 sg13g2_o21ai_1 _5312_ (.B1(_0987_),
    .Y(_0993_),
    .A1(_0982_),
    .A2(_0988_));
 sg13g2_o21ai_1 _5313_ (.B1(_0882_),
    .Y(_0994_),
    .A1(_0973_),
    .A2(_0975_));
 sg13g2_a221oi_1 _5314_ (.B2(_0977_),
    .C1(_0994_),
    .B1(_0993_),
    .A1(_0964_),
    .Y(_0995_),
    .A2(_0992_));
 sg13g2_nor3_1 _5315_ (.A(net298),
    .B(net1209),
    .C(_0995_),
    .Y(_0107_));
 sg13g2_and2_1 _5316_ (.A(net1337),
    .B(net302),
    .X(_0108_));
 sg13g2_o21ai_1 _5317_ (.B1(net1106),
    .Y(_0996_),
    .A1(net1092),
    .A2(net1229));
 sg13g2_nor2b_1 _5318_ (.A(net1229),
    .B_N(net1098),
    .Y(_0997_));
 sg13g2_nor2_1 _5319_ (.A(_0996_),
    .B(_0997_),
    .Y(_0998_));
 sg13g2_inv_1 _5320_ (.Y(_0999_),
    .A(_0998_));
 sg13g2_o21ai_1 _5321_ (.B1(_0999_),
    .Y(_1000_),
    .A1(net1105),
    .A2(_0879_));
 sg13g2_or2_1 _5322_ (.X(_1001_),
    .B(net1098),
    .A(\s0.was_valid_out[11] [0]));
 sg13g2_o21ai_1 _5323_ (.B1(net938),
    .Y(_1002_),
    .A1(\s0.was_valid_out[11] [0]),
    .A2(net1110));
 sg13g2_o21ai_1 _5324_ (.B1(_1002_),
    .Y(_1003_),
    .A1(net1092),
    .A2(_0996_));
 sg13g2_a21oi_1 _5325_ (.A1(_0998_),
    .A2(_1001_),
    .Y(_1004_),
    .B1(_1003_));
 sg13g2_o21ai_1 _5326_ (.B1(net1336),
    .Y(_1005_),
    .A1(net408),
    .A2(_1000_));
 sg13g2_nor2_1 _5327_ (.A(_1004_),
    .B(_1005_),
    .Y(_0109_));
 sg13g2_nor2_1 _5328_ (.A(net1220),
    .B(_1000_),
    .Y(_0110_));
 sg13g2_mux2_1 _5329_ (.A0(\s0.data_out[11][0] ),
    .A1(\s0.data_out[12][0] ),
    .S(net1108),
    .X(_1006_));
 sg13g2_nand2_1 _5330_ (.Y(_1007_),
    .A(net938),
    .B(_1006_));
 sg13g2_and2_1 _5331_ (.A(net1088),
    .B(\s0.data_out[11][0] ),
    .X(_1008_));
 sg13g2_nor2b_1 _5332_ (.A(net1088),
    .B_N(net1074),
    .Y(_1009_));
 sg13g2_o21ai_1 _5333_ (.B1(net1102),
    .Y(_1010_),
    .A1(_1008_),
    .A2(_1009_));
 sg13g2_nand3_1 _5334_ (.B(_1007_),
    .C(_1010_),
    .A(net1335),
    .Y(_1011_));
 sg13g2_o21ai_1 _5335_ (.B1(_1011_),
    .Y(_1012_),
    .A1(net1335),
    .A2(net473));
 sg13g2_inv_1 _5336_ (.Y(_0111_),
    .A(_1012_));
 sg13g2_nand2b_1 _5337_ (.Y(_1013_),
    .B(\s0.data_out[11][1] ),
    .A_N(net1109));
 sg13g2_a21oi_1 _5338_ (.A1(_0948_),
    .A2(_1013_),
    .Y(_1014_),
    .B1(net1102));
 sg13g2_nor2b_1 _5339_ (.A(net1088),
    .B_N(net1070),
    .Y(_1015_));
 sg13g2_a21oi_1 _5340_ (.A1(net1088),
    .A2(\s0.data_out[11][1] ),
    .Y(_1016_),
    .B1(_1015_));
 sg13g2_o21ai_1 _5341_ (.B1(net1334),
    .Y(_1017_),
    .A1(net938),
    .A2(_1016_));
 sg13g2_or2_1 _5342_ (.X(_1018_),
    .B(net528),
    .A(net1334));
 sg13g2_o21ai_1 _5343_ (.B1(_1018_),
    .Y(_1019_),
    .A1(_1014_),
    .A2(_1017_));
 sg13g2_inv_1 _5344_ (.Y(_0112_),
    .A(net529));
 sg13g2_nand2b_1 _5345_ (.Y(_1020_),
    .B(\s0.data_out[11][2] ),
    .A_N(net1109));
 sg13g2_a21oi_1 _5346_ (.A1(_0944_),
    .A2(_1020_),
    .Y(_1021_),
    .B1(net1102));
 sg13g2_nor2b_1 _5347_ (.A(net1089),
    .B_N(net1066),
    .Y(_1022_));
 sg13g2_a21oi_1 _5348_ (.A1(net1088),
    .A2(\s0.data_out[11][2] ),
    .Y(_1023_),
    .B1(_1022_));
 sg13g2_o21ai_1 _5349_ (.B1(net1334),
    .Y(_1024_),
    .A1(net938),
    .A2(_1023_));
 sg13g2_or2_1 _5350_ (.X(_1025_),
    .B(net504),
    .A(net1332));
 sg13g2_o21ai_1 _5351_ (.B1(_1025_),
    .Y(_1026_),
    .A1(_1021_),
    .A2(_1024_));
 sg13g2_inv_1 _5352_ (.Y(_0113_),
    .A(net505));
 sg13g2_mux2_1 _5353_ (.A0(\s0.data_out[11][3] ),
    .A1(\s0.data_out[12][3] ),
    .S(net1108),
    .X(_1027_));
 sg13g2_nand2_1 _5354_ (.Y(_1028_),
    .A(net938),
    .B(_1027_));
 sg13g2_and2_1 _5355_ (.A(net1088),
    .B(net613),
    .X(_1029_));
 sg13g2_nor2b_1 _5356_ (.A(net1089),
    .B_N(net1062),
    .Y(_1030_));
 sg13g2_o21ai_1 _5357_ (.B1(net1103),
    .Y(_1031_),
    .A1(_1029_),
    .A2(_1030_));
 sg13g2_nand3_1 _5358_ (.B(_1028_),
    .C(_1031_),
    .A(net1334),
    .Y(_1032_));
 sg13g2_o21ai_1 _5359_ (.B1(net614),
    .Y(_1033_),
    .A1(net1334),
    .A2(net472));
 sg13g2_inv_1 _5360_ (.Y(_0114_),
    .A(_1033_));
 sg13g2_nand2b_1 _5361_ (.Y(_1034_),
    .B(net330),
    .A_N(net1110));
 sg13g2_a21oi_1 _5362_ (.A1(_0978_),
    .A2(_1034_),
    .Y(_1035_),
    .B1(net1103));
 sg13g2_nor2b_1 _5363_ (.A(net1092),
    .B_N(net1059),
    .Y(_1036_));
 sg13g2_a21oi_1 _5364_ (.A1(net1092),
    .A2(net330),
    .Y(_1037_),
    .B1(_1036_));
 sg13g2_o21ai_1 _5365_ (.B1(net1337),
    .Y(_1038_),
    .A1(net938),
    .A2(_1037_));
 sg13g2_or2_1 _5366_ (.X(_1039_),
    .B(net556),
    .A(net1337));
 sg13g2_o21ai_1 _5367_ (.B1(_1039_),
    .Y(_1040_),
    .A1(net331),
    .A2(_1038_));
 sg13g2_inv_1 _5368_ (.Y(_0115_),
    .A(_1040_));
 sg13g2_nand2b_1 _5369_ (.Y(_1041_),
    .B(\s0.data_out[11][5] ),
    .A_N(net1110));
 sg13g2_a21oi_1 _5370_ (.A1(_0983_),
    .A2(_1041_),
    .Y(_1042_),
    .B1(net1105));
 sg13g2_nor2b_1 _5371_ (.A(net1092),
    .B_N(net1055),
    .Y(_1043_));
 sg13g2_a21oi_1 _5372_ (.A1(net1091),
    .A2(\s0.data_out[11][5] ),
    .Y(_1044_),
    .B1(_1043_));
 sg13g2_o21ai_1 _5373_ (.B1(net1339),
    .Y(_1045_),
    .A1(net938),
    .A2(_1044_));
 sg13g2_or2_1 _5374_ (.X(_1046_),
    .B(net501),
    .A(net1336));
 sg13g2_o21ai_1 _5375_ (.B1(_1046_),
    .Y(_1047_),
    .A1(_1042_),
    .A2(_1045_));
 sg13g2_inv_1 _5376_ (.Y(_0116_),
    .A(net502));
 sg13g2_nand2b_1 _5377_ (.Y(_1048_),
    .B(net527),
    .A_N(net1110));
 sg13g2_a21oi_1 _5378_ (.A1(_0969_),
    .A2(_1048_),
    .Y(_1049_),
    .B1(net1105));
 sg13g2_nor2b_1 _5379_ (.A(net1091),
    .B_N(net1051),
    .Y(_1050_));
 sg13g2_a21oi_1 _5380_ (.A1(net1091),
    .A2(net527),
    .Y(_1051_),
    .B1(_1050_));
 sg13g2_o21ai_1 _5381_ (.B1(net1336),
    .Y(_1052_),
    .A1(net938),
    .A2(_1051_));
 sg13g2_or2_1 _5382_ (.X(_1053_),
    .B(net588),
    .A(net1336));
 sg13g2_o21ai_1 _5383_ (.B1(_1053_),
    .Y(_1054_),
    .A1(_1049_),
    .A2(_1052_));
 sg13g2_inv_1 _5384_ (.Y(_0117_),
    .A(_1054_));
 sg13g2_nand2b_1 _5385_ (.Y(_1055_),
    .B(net540),
    .A_N(net1110));
 sg13g2_a21oi_1 _5386_ (.A1(_0965_),
    .A2(_1055_),
    .Y(_1056_),
    .B1(net1105));
 sg13g2_nor2b_1 _5387_ (.A(net1091),
    .B_N(net1047),
    .Y(_1057_));
 sg13g2_a21oi_1 _5388_ (.A1(net1091),
    .A2(net540),
    .Y(_1058_),
    .B1(_1057_));
 sg13g2_o21ai_1 _5389_ (.B1(net1336),
    .Y(_1059_),
    .A1(_2451_),
    .A2(_1058_));
 sg13g2_or2_1 _5390_ (.X(_1060_),
    .B(net594),
    .A(net1336));
 sg13g2_o21ai_1 _5391_ (.B1(_1060_),
    .Y(_1061_),
    .A1(_1056_),
    .A2(_1059_));
 sg13g2_inv_1 _5392_ (.Y(_0118_),
    .A(_1061_));
 sg13g2_nand2_1 _5393_ (.Y(_1062_),
    .A(net1099),
    .B(net568));
 sg13g2_mux2_1 _5394_ (.A0(\s0.data_out[12][2] ),
    .A1(\s0.data_out[11][2] ),
    .S(net1096),
    .X(_1063_));
 sg13g2_a21o_1 _5395_ (.A2(_1063_),
    .A1(net1089),
    .B1(_1022_),
    .X(_1064_));
 sg13g2_a21oi_1 _5396_ (.A1(net1103),
    .A2(_1064_),
    .Y(_1065_),
    .B1(_1021_));
 sg13g2_nor2_1 _5397_ (.A(net1270),
    .B(_1065_),
    .Y(_1066_));
 sg13g2_nand2_1 _5398_ (.Y(_1067_),
    .A(net1099),
    .B(net536));
 sg13g2_mux2_1 _5399_ (.A0(\s0.data_out[12][1] ),
    .A1(\s0.data_out[11][1] ),
    .S(net1096),
    .X(_1068_));
 sg13g2_a21o_1 _5400_ (.A2(_1068_),
    .A1(net1088),
    .B1(_1015_),
    .X(_1069_));
 sg13g2_a21oi_1 _5401_ (.A1(net1102),
    .A2(_1069_),
    .Y(_1070_),
    .B1(_1014_));
 sg13g2_mux2_1 _5402_ (.A0(\s0.data_out[12][0] ),
    .A1(\s0.data_out[11][0] ),
    .S(net1096),
    .X(_1071_));
 sg13g2_a21oi_1 _5403_ (.A1(net1088),
    .A2(_1071_),
    .Y(_1072_),
    .B1(_1009_));
 sg13g2_nand2b_1 _5404_ (.Y(_1073_),
    .B(net1102),
    .A_N(_1072_));
 sg13g2_nor2_1 _5405_ (.A(net1279),
    .B(_1070_),
    .Y(_1074_));
 sg13g2_a221oi_1 _5406_ (.B2(_1007_),
    .C1(net1282),
    .B1(_1073_),
    .A1(net1279),
    .Y(_1075_),
    .A2(_1070_));
 sg13g2_nor3_1 _5407_ (.A(_1066_),
    .B(_1074_),
    .C(_1075_),
    .Y(_1076_));
 sg13g2_nand2_1 _5408_ (.Y(_1077_),
    .A(net1096),
    .B(net486));
 sg13g2_o21ai_1 _5409_ (.B1(_1077_),
    .Y(_1078_),
    .A1(net1096),
    .A2(_2488_));
 sg13g2_a21oi_1 _5410_ (.A1(net1089),
    .A2(_1078_),
    .Y(_1079_),
    .B1(_1030_));
 sg13g2_nand2b_1 _5411_ (.Y(_1080_),
    .B(net1103),
    .A_N(_1079_));
 sg13g2_and2_1 _5412_ (.A(_1028_),
    .B(_1080_),
    .X(_1081_));
 sg13g2_a221oi_1 _5413_ (.B2(net1265),
    .C1(_1076_),
    .B1(_1081_),
    .A1(net1270),
    .Y(_1082_),
    .A2(_1065_));
 sg13g2_nand2_1 _5414_ (.Y(_1083_),
    .A(net1097),
    .B(net540));
 sg13g2_mux2_1 _5415_ (.A0(\s0.data_out[12][7] ),
    .A1(\s0.data_out[11][7] ),
    .S(net1098),
    .X(_1084_));
 sg13g2_a21o_1 _5416_ (.A2(_1084_),
    .A1(net1091),
    .B1(_1057_),
    .X(_1085_));
 sg13g2_a21oi_1 _5417_ (.A1(net1105),
    .A2(_1085_),
    .Y(_1086_),
    .B1(_1056_));
 sg13g2_nand2_1 _5418_ (.Y(_1087_),
    .A(net1097),
    .B(net527));
 sg13g2_mux2_1 _5419_ (.A0(\s0.data_out[12][6] ),
    .A1(\s0.data_out[11][6] ),
    .S(net1098),
    .X(_1088_));
 sg13g2_a21o_1 _5420_ (.A2(_1088_),
    .A1(net1091),
    .B1(_1050_),
    .X(_1089_));
 sg13g2_a21oi_1 _5421_ (.A1(net1105),
    .A2(_1089_),
    .Y(_1090_),
    .B1(_1049_));
 sg13g2_a22oi_1 _5422_ (.Y(_1091_),
    .B1(_1090_),
    .B2(net1242),
    .A2(_1086_),
    .A1(net1236));
 sg13g2_or2_1 _5423_ (.X(_1092_),
    .B(_1086_),
    .A(net1236));
 sg13g2_nor2_1 _5424_ (.A(net1242),
    .B(_1090_),
    .Y(_1093_));
 sg13g2_nand3b_1 _5425_ (.B(_1091_),
    .C(_1092_),
    .Y(_1094_),
    .A_N(_1093_));
 sg13g2_nand2_1 _5426_ (.Y(_1095_),
    .A(net1097),
    .B(net330));
 sg13g2_mux2_1 _5427_ (.A0(\s0.data_out[12][4] ),
    .A1(\s0.data_out[11][4] ),
    .S(net1098),
    .X(_1096_));
 sg13g2_a21o_1 _5428_ (.A2(_1096_),
    .A1(net1092),
    .B1(_1036_),
    .X(_1097_));
 sg13g2_a21oi_1 _5429_ (.A1(net1103),
    .A2(_1097_),
    .Y(_1098_),
    .B1(_1035_));
 sg13g2_nand2_1 _5430_ (.Y(_1099_),
    .A(net1256),
    .B(_1098_));
 sg13g2_nand2_1 _5431_ (.Y(_1100_),
    .A(net1098),
    .B(net541));
 sg13g2_mux2_1 _5432_ (.A0(\s0.data_out[12][5] ),
    .A1(\s0.data_out[11][5] ),
    .S(net1098),
    .X(_1101_));
 sg13g2_a21o_1 _5433_ (.A2(_1101_),
    .A1(net1091),
    .B1(_1043_),
    .X(_1102_));
 sg13g2_a21oi_1 _5434_ (.A1(net1105),
    .A2(_1102_),
    .Y(_1103_),
    .B1(_1042_));
 sg13g2_nand2_1 _5435_ (.Y(_1104_),
    .A(net1251),
    .B(_1103_));
 sg13g2_or2_1 _5436_ (.X(_1105_),
    .B(_1103_),
    .A(net1251));
 sg13g2_or2_1 _5437_ (.X(_1106_),
    .B(_1098_),
    .A(net1256));
 sg13g2_o21ai_1 _5438_ (.B1(_1099_),
    .Y(_1107_),
    .A1(net1265),
    .A2(_1081_));
 sg13g2_nand3_1 _5439_ (.B(_1105_),
    .C(_1106_),
    .A(_1104_),
    .Y(_1108_));
 sg13g2_or4_1 _5440_ (.A(_1082_),
    .B(_1094_),
    .C(_1107_),
    .D(_1108_),
    .X(_1109_));
 sg13g2_nand2b_1 _5441_ (.Y(_1110_),
    .B(_1105_),
    .A_N(_1099_));
 sg13g2_a21oi_1 _5442_ (.A1(_1104_),
    .A2(_1110_),
    .Y(_1111_),
    .B1(_1094_));
 sg13g2_nor2b_1 _5443_ (.A(_1091_),
    .B_N(_1092_),
    .Y(_1112_));
 sg13g2_nor3_1 _5444_ (.A(_1000_),
    .B(_1111_),
    .C(_1112_),
    .Y(_1113_));
 sg13g2_or2_1 _5445_ (.X(_1114_),
    .B(net1209),
    .A(net302));
 sg13g2_a21oi_1 _5446_ (.A1(_1109_),
    .A2(_1113_),
    .Y(_0119_),
    .B1(_1114_));
 sg13g2_and2_1 _5447_ (.A(net316),
    .B(net1345),
    .X(_0120_));
 sg13g2_o21ai_1 _5448_ (.B1(net1093),
    .Y(_1115_),
    .A1(net1229),
    .A2(net1080));
 sg13g2_nor2b_1 _5449_ (.A(net1229),
    .B_N(net1085),
    .Y(_1116_));
 sg13g2_nor2_1 _5450_ (.A(_1115_),
    .B(_1116_),
    .Y(_1117_));
 sg13g2_nor2_1 _5451_ (.A(net1094),
    .B(_0997_),
    .Y(_1118_));
 sg13g2_or2_1 _5452_ (.X(_1119_),
    .B(_1118_),
    .A(_1117_));
 sg13g2_or2_1 _5453_ (.X(_1120_),
    .B(net1085),
    .A(net379));
 sg13g2_o21ai_1 _5454_ (.B1(net939),
    .Y(_1121_),
    .A1(net379),
    .A2(net1097));
 sg13g2_o21ai_1 _5455_ (.B1(_1121_),
    .Y(_1122_),
    .A1(net1080),
    .A2(_1115_));
 sg13g2_a21oi_1 _5456_ (.A1(_1117_),
    .A2(_1120_),
    .Y(_1123_),
    .B1(_1122_));
 sg13g2_o21ai_1 _5457_ (.B1(net1336),
    .Y(_1124_),
    .A1(net413),
    .A2(_1119_));
 sg13g2_nor2_1 _5458_ (.A(_1123_),
    .B(_1124_),
    .Y(_0121_));
 sg13g2_nor2_1 _5459_ (.A(net1221),
    .B(_1119_),
    .Y(_0122_));
 sg13g2_mux2_1 _5460_ (.A0(\s0.data_out[10][0] ),
    .A1(\s0.data_out[11][0] ),
    .S(net1096),
    .X(_1125_));
 sg13g2_nand2_1 _5461_ (.Y(_1126_),
    .A(net939),
    .B(_1125_));
 sg13g2_and2_1 _5462_ (.A(net1077),
    .B(\s0.data_out[10][0] ),
    .X(_1127_));
 sg13g2_nor2b_1 _5463_ (.A(net1077),
    .B_N(net1074),
    .Y(_1128_));
 sg13g2_o21ai_1 _5464_ (.B1(net1090),
    .Y(_1129_),
    .A1(_1127_),
    .A2(_1128_));
 sg13g2_nand3_1 _5465_ (.B(_1126_),
    .C(_1129_),
    .A(net1335),
    .Y(_1130_));
 sg13g2_o21ai_1 _5466_ (.B1(_1130_),
    .Y(_1131_),
    .A1(net1335),
    .A2(net452));
 sg13g2_inv_1 _5467_ (.Y(_0123_),
    .A(_1131_));
 sg13g2_nand2b_1 _5468_ (.Y(_1132_),
    .B(net418),
    .A_N(net1099));
 sg13g2_a21oi_1 _5469_ (.A1(_1067_),
    .A2(_1132_),
    .Y(_1133_),
    .B1(net1090));
 sg13g2_nor2b_1 _5470_ (.A(net1077),
    .B_N(net1070),
    .Y(_1134_));
 sg13g2_a21oi_1 _5471_ (.A1(net1077),
    .A2(net418),
    .Y(_1135_),
    .B1(_1134_));
 sg13g2_o21ai_1 _5472_ (.B1(net1335),
    .Y(_1136_),
    .A1(net939),
    .A2(_1135_));
 sg13g2_or2_1 _5473_ (.X(_1137_),
    .B(net536),
    .A(net1334));
 sg13g2_o21ai_1 _5474_ (.B1(_1137_),
    .Y(_1138_),
    .A1(_1133_),
    .A2(_1136_));
 sg13g2_inv_1 _5475_ (.Y(_0124_),
    .A(_1138_));
 sg13g2_nand2b_1 _5476_ (.Y(_1139_),
    .B(net506),
    .A_N(net1096));
 sg13g2_a21oi_1 _5477_ (.A1(_1062_),
    .A2(_1139_),
    .Y(_1140_),
    .B1(net1090));
 sg13g2_nor2b_1 _5478_ (.A(net1079),
    .B_N(net1067),
    .Y(_1141_));
 sg13g2_a21oi_1 _5479_ (.A1(net1078),
    .A2(net506),
    .Y(_1142_),
    .B1(_1141_));
 sg13g2_o21ai_1 _5480_ (.B1(net1344),
    .Y(_1143_),
    .A1(net939),
    .A2(_1142_));
 sg13g2_or2_1 _5481_ (.X(_1144_),
    .B(net568),
    .A(net1337));
 sg13g2_o21ai_1 _5482_ (.B1(_1144_),
    .Y(_1145_),
    .A1(_1140_),
    .A2(_1143_));
 sg13g2_inv_1 _5483_ (.Y(_0125_),
    .A(_1145_));
 sg13g2_nand2b_1 _5484_ (.Y(_1146_),
    .B(net436),
    .A_N(net1096));
 sg13g2_a21oi_1 _5485_ (.A1(_1077_),
    .A2(_1146_),
    .Y(_1147_),
    .B1(net1090));
 sg13g2_nor2b_1 _5486_ (.A(net1079),
    .B_N(net1062),
    .Y(_1148_));
 sg13g2_a21oi_1 _5487_ (.A1(net1078),
    .A2(net436),
    .Y(_1149_),
    .B1(_1148_));
 sg13g2_o21ai_1 _5488_ (.B1(net1335),
    .Y(_1150_),
    .A1(net939),
    .A2(_1149_));
 sg13g2_or2_1 _5489_ (.X(_1151_),
    .B(net486),
    .A(net1335));
 sg13g2_o21ai_1 _5490_ (.B1(_1151_),
    .Y(_1152_),
    .A1(_1147_),
    .A2(_1150_));
 sg13g2_inv_1 _5491_ (.Y(_0126_),
    .A(_1152_));
 sg13g2_nand2b_1 _5492_ (.Y(_1153_),
    .B(net429),
    .A_N(net1097));
 sg13g2_a21oi_1 _5493_ (.A1(_1095_),
    .A2(_1153_),
    .Y(_1154_),
    .B1(net1093));
 sg13g2_nor2b_1 _5494_ (.A(net1081),
    .B_N(net1059),
    .Y(_1155_));
 sg13g2_a21oi_1 _5495_ (.A1(net1081),
    .A2(net429),
    .Y(_1156_),
    .B1(_1155_));
 sg13g2_o21ai_1 _5496_ (.B1(net1337),
    .Y(_1157_),
    .A1(net939),
    .A2(_1156_));
 sg13g2_or2_1 _5497_ (.X(_1158_),
    .B(net330),
    .A(net1337));
 sg13g2_o21ai_1 _5498_ (.B1(_1158_),
    .Y(_1159_),
    .A1(_1154_),
    .A2(_1157_));
 sg13g2_inv_1 _5499_ (.Y(_0127_),
    .A(_1159_));
 sg13g2_nand2b_1 _5500_ (.Y(_1160_),
    .B(net481),
    .A_N(net1097));
 sg13g2_a21oi_1 _5501_ (.A1(_1100_),
    .A2(_1160_),
    .Y(_1161_),
    .B1(net1093));
 sg13g2_nor2b_1 _5502_ (.A(net1080),
    .B_N(net1055),
    .Y(_1162_));
 sg13g2_a21oi_1 _5503_ (.A1(net1080),
    .A2(net481),
    .Y(_1163_),
    .B1(_1162_));
 sg13g2_o21ai_1 _5504_ (.B1(net1345),
    .Y(_1164_),
    .A1(net939),
    .A2(_1163_));
 sg13g2_or2_1 _5505_ (.X(_1165_),
    .B(net541),
    .A(net1336));
 sg13g2_o21ai_1 _5506_ (.B1(_1165_),
    .Y(_1166_),
    .A1(_1161_),
    .A2(_1164_));
 sg13g2_inv_1 _5507_ (.Y(_0128_),
    .A(_1166_));
 sg13g2_nand2b_1 _5508_ (.Y(_1167_),
    .B(net521),
    .A_N(net1097));
 sg13g2_a21oi_1 _5509_ (.A1(_1087_),
    .A2(_1167_),
    .Y(_1168_),
    .B1(net1093));
 sg13g2_nor2b_1 _5510_ (.A(net1081),
    .B_N(net1051),
    .Y(_1169_));
 sg13g2_a21oi_1 _5511_ (.A1(net1081),
    .A2(net521),
    .Y(_1170_),
    .B1(_1169_));
 sg13g2_o21ai_1 _5512_ (.B1(net1344),
    .Y(_1171_),
    .A1(net939),
    .A2(_1170_));
 sg13g2_or2_1 _5513_ (.X(_1172_),
    .B(net527),
    .A(net1345));
 sg13g2_o21ai_1 _5514_ (.B1(_1172_),
    .Y(_1173_),
    .A1(_1168_),
    .A2(_1171_));
 sg13g2_inv_1 _5515_ (.Y(_0129_),
    .A(_1173_));
 sg13g2_nand2b_1 _5516_ (.Y(_1174_),
    .B(net531),
    .A_N(net1097));
 sg13g2_a21oi_1 _5517_ (.A1(_1083_),
    .A2(_1174_),
    .Y(_1175_),
    .B1(net1093));
 sg13g2_nor2b_1 _5518_ (.A(net1080),
    .B_N(net1047),
    .Y(_1176_));
 sg13g2_a21oi_1 _5519_ (.A1(net1080),
    .A2(net531),
    .Y(_1177_),
    .B1(_1176_));
 sg13g2_o21ai_1 _5520_ (.B1(net1344),
    .Y(_1178_),
    .A1(_2448_),
    .A2(_1177_));
 sg13g2_or2_1 _5521_ (.X(_1179_),
    .B(net540),
    .A(net1345));
 sg13g2_o21ai_1 _5522_ (.B1(_1179_),
    .Y(_1180_),
    .A1(_1175_),
    .A2(_1178_));
 sg13g2_inv_1 _5523_ (.Y(_0130_),
    .A(_1180_));
 sg13g2_nand2_1 _5524_ (.Y(_1181_),
    .A(net1084),
    .B(net506));
 sg13g2_mux2_1 _5525_ (.A0(\s0.data_out[11][2] ),
    .A1(\s0.data_out[10][2] ),
    .S(net1084),
    .X(_1182_));
 sg13g2_a21o_1 _5526_ (.A2(_1182_),
    .A1(net1078),
    .B1(_1141_),
    .X(_1183_));
 sg13g2_a21oi_1 _5527_ (.A1(net1095),
    .A2(_1183_),
    .Y(_1184_),
    .B1(_1140_));
 sg13g2_nor2_1 _5528_ (.A(net1270),
    .B(_1184_),
    .Y(_1185_));
 sg13g2_mux2_1 _5529_ (.A0(\s0.data_out[11][1] ),
    .A1(\s0.data_out[10][1] ),
    .S(net1084),
    .X(_1186_));
 sg13g2_a21o_1 _5530_ (.A2(_1186_),
    .A1(net1077),
    .B1(_1134_),
    .X(_1187_));
 sg13g2_a21oi_1 _5531_ (.A1(net1090),
    .A2(_1187_),
    .Y(_1188_),
    .B1(_1133_));
 sg13g2_mux2_1 _5532_ (.A0(\s0.data_out[11][0] ),
    .A1(\s0.data_out[10][0] ),
    .S(net1084),
    .X(_1189_));
 sg13g2_a21oi_1 _5533_ (.A1(net1077),
    .A2(_1189_),
    .Y(_1190_),
    .B1(_1128_));
 sg13g2_nand2b_1 _5534_ (.Y(_1191_),
    .B(net1090),
    .A_N(_1190_));
 sg13g2_nor2_1 _5535_ (.A(net1278),
    .B(_1188_),
    .Y(_1192_));
 sg13g2_a221oi_1 _5536_ (.B2(_1126_),
    .C1(net1283),
    .B1(_1191_),
    .A1(net1278),
    .Y(_1193_),
    .A2(_1188_));
 sg13g2_nor3_1 _5537_ (.A(_1185_),
    .B(_1192_),
    .C(_1193_),
    .Y(_1194_));
 sg13g2_mux2_1 _5538_ (.A0(\s0.data_out[11][3] ),
    .A1(\s0.data_out[10][3] ),
    .S(net1084),
    .X(_1195_));
 sg13g2_a21o_1 _5539_ (.A2(_1195_),
    .A1(net1078),
    .B1(_1148_),
    .X(_1196_));
 sg13g2_a21oi_1 _5540_ (.A1(net1095),
    .A2(_1196_),
    .Y(_1197_),
    .B1(_1147_));
 sg13g2_a221oi_1 _5541_ (.B2(net1266),
    .C1(_1194_),
    .B1(_1197_),
    .A1(net1270),
    .Y(_1198_),
    .A2(_1184_));
 sg13g2_nand2_1 _5542_ (.Y(_1199_),
    .A(net1085),
    .B(net531));
 sg13g2_mux2_1 _5543_ (.A0(\s0.data_out[11][7] ),
    .A1(\s0.data_out[10][7] ),
    .S(net1085),
    .X(_1200_));
 sg13g2_a21o_1 _5544_ (.A2(_1200_),
    .A1(net1080),
    .B1(_1176_),
    .X(_1201_));
 sg13g2_a21oi_1 _5545_ (.A1(net1094),
    .A2(_1201_),
    .Y(_1202_),
    .B1(_1175_));
 sg13g2_nand2_1 _5546_ (.Y(_1203_),
    .A(net1086),
    .B(net521));
 sg13g2_mux2_1 _5547_ (.A0(\s0.data_out[11][6] ),
    .A1(\s0.data_out[10][6] ),
    .S(net1085),
    .X(_1204_));
 sg13g2_a21o_1 _5548_ (.A2(_1204_),
    .A1(net1081),
    .B1(_1169_),
    .X(_1205_));
 sg13g2_a21oi_1 _5549_ (.A1(net1094),
    .A2(_1205_),
    .Y(_1206_),
    .B1(_1168_));
 sg13g2_a22oi_1 _5550_ (.Y(_1207_),
    .B1(_1206_),
    .B2(net1242),
    .A2(_1202_),
    .A1(net1236));
 sg13g2_or2_1 _5551_ (.X(_1208_),
    .B(_1206_),
    .A(net1243));
 sg13g2_or2_1 _5552_ (.X(_1209_),
    .B(_1202_),
    .A(net1237));
 sg13g2_nand3_1 _5553_ (.B(_1208_),
    .C(_1209_),
    .A(_1207_),
    .Y(_1210_));
 sg13g2_mux2_1 _5554_ (.A0(\s0.data_out[11][4] ),
    .A1(\s0.data_out[10][4] ),
    .S(net1085),
    .X(_1211_));
 sg13g2_a21o_1 _5555_ (.A2(_1211_),
    .A1(net1081),
    .B1(_1155_),
    .X(_1212_));
 sg13g2_a21oi_1 _5556_ (.A1(net1093),
    .A2(_1212_),
    .Y(_1213_),
    .B1(_1154_));
 sg13g2_nand2_1 _5557_ (.Y(_1214_),
    .A(net1086),
    .B(\s0.data_out[10][5] ));
 sg13g2_mux2_1 _5558_ (.A0(\s0.data_out[11][5] ),
    .A1(\s0.data_out[10][5] ),
    .S(net1085),
    .X(_1215_));
 sg13g2_a21o_1 _5559_ (.A2(_1215_),
    .A1(net1080),
    .B1(_1162_),
    .X(_1216_));
 sg13g2_a21oi_1 _5560_ (.A1(net1093),
    .A2(_1216_),
    .Y(_1217_),
    .B1(_1161_));
 sg13g2_a22oi_1 _5561_ (.Y(_1218_),
    .B1(_1217_),
    .B2(net1252),
    .A2(_1213_),
    .A1(net1256));
 sg13g2_nor2_1 _5562_ (.A(net1256),
    .B(_1213_),
    .Y(_1219_));
 sg13g2_nor2_1 _5563_ (.A(net1252),
    .B(_1217_),
    .Y(_1220_));
 sg13g2_nor2_1 _5564_ (.A(net1265),
    .B(_1197_),
    .Y(_1221_));
 sg13g2_nor3_1 _5565_ (.A(_1219_),
    .B(_1220_),
    .C(_1221_),
    .Y(_1222_));
 sg13g2_nand2_1 _5566_ (.Y(_1223_),
    .A(_1218_),
    .B(_1222_));
 sg13g2_or3_1 _5567_ (.A(_1198_),
    .B(_1210_),
    .C(_1223_),
    .X(_1224_));
 sg13g2_nor3_1 _5568_ (.A(_1210_),
    .B(_1218_),
    .C(_1220_),
    .Y(_1225_));
 sg13g2_nor2b_1 _5569_ (.A(_1207_),
    .B_N(_1209_),
    .Y(_1226_));
 sg13g2_nor3_1 _5570_ (.A(_1119_),
    .B(_1225_),
    .C(_1226_),
    .Y(_1227_));
 sg13g2_or2_1 _5571_ (.X(_1228_),
    .B(net1210),
    .A(net316));
 sg13g2_a21oi_1 _5572_ (.A1(_1224_),
    .A2(_1227_),
    .Y(_0131_),
    .B1(_1228_));
 sg13g2_and2_1 _5573_ (.A(net1346),
    .B(net315),
    .X(_0132_));
 sg13g2_o21ai_1 _5574_ (.B1(net1082),
    .Y(_1229_),
    .A1(net1229),
    .A2(net1039));
 sg13g2_nor2b_1 _5575_ (.A(net1229),
    .B_N(net1044),
    .Y(_1230_));
 sg13g2_nor2_1 _5576_ (.A(_1229_),
    .B(_1230_),
    .Y(_1231_));
 sg13g2_inv_1 _5577_ (.Y(_1232_),
    .A(_1231_));
 sg13g2_o21ai_1 _5578_ (.B1(_1232_),
    .Y(_1233_),
    .A1(net1082),
    .A2(_1116_));
 sg13g2_or2_1 _5579_ (.X(_1234_),
    .B(net1043),
    .A(\s0.was_valid_out[9] [0]));
 sg13g2_o21ai_1 _5580_ (.B1(net934),
    .Y(_1235_),
    .A1(\s0.was_valid_out[9] [0]),
    .A2(net1085));
 sg13g2_o21ai_1 _5581_ (.B1(_1235_),
    .Y(_1236_),
    .A1(net1038),
    .A2(_1229_));
 sg13g2_a21oi_1 _5582_ (.A1(_1231_),
    .A2(_1234_),
    .Y(_1237_),
    .B1(_1236_));
 sg13g2_o21ai_1 _5583_ (.B1(net1344),
    .Y(_1238_),
    .A1(net379),
    .A2(_1233_));
 sg13g2_nor2_1 _5584_ (.A(_1237_),
    .B(_1238_),
    .Y(_0133_));
 sg13g2_nor2_1 _5585_ (.A(net1221),
    .B(_1233_),
    .Y(_0134_));
 sg13g2_mux2_1 _5586_ (.A0(\s0.data_out[9][0] ),
    .A1(\s0.data_out[10][0] ),
    .S(net1084),
    .X(_1239_));
 sg13g2_nand2_1 _5587_ (.Y(_1240_),
    .A(net934),
    .B(_1239_));
 sg13g2_and2_1 _5588_ (.A(net1035),
    .B(\s0.data_out[9][0] ),
    .X(_1241_));
 sg13g2_nor2b_1 _5589_ (.A(net1035),
    .B_N(net1074),
    .Y(_1242_));
 sg13g2_o21ai_1 _5590_ (.B1(net1077),
    .Y(_1243_),
    .A1(_1241_),
    .A2(_1242_));
 sg13g2_nand3_1 _5591_ (.B(_1240_),
    .C(_1243_),
    .A(net1340),
    .Y(_1244_));
 sg13g2_o21ai_1 _5592_ (.B1(_1244_),
    .Y(_1245_),
    .A1(net1340),
    .A2(net404));
 sg13g2_inv_1 _5593_ (.Y(_0135_),
    .A(_1245_));
 sg13g2_mux2_1 _5594_ (.A0(\s0.data_out[9][1] ),
    .A1(\s0.data_out[10][1] ),
    .S(net1084),
    .X(_1246_));
 sg13g2_nand2_1 _5595_ (.Y(_1247_),
    .A(net934),
    .B(_1246_));
 sg13g2_and2_1 _5596_ (.A(net1036),
    .B(\s0.data_out[9][1] ),
    .X(_1248_));
 sg13g2_nor2b_1 _5597_ (.A(net1036),
    .B_N(net1071),
    .Y(_1249_));
 sg13g2_o21ai_1 _5598_ (.B1(net1077),
    .Y(_1250_),
    .A1(_1248_),
    .A2(_1249_));
 sg13g2_nand3_1 _5599_ (.B(_1247_),
    .C(_1250_),
    .A(net1341),
    .Y(_1251_));
 sg13g2_o21ai_1 _5600_ (.B1(_1251_),
    .Y(_1252_),
    .A1(net1341),
    .A2(net418));
 sg13g2_inv_1 _5601_ (.Y(_0136_),
    .A(_1252_));
 sg13g2_nand2b_1 _5602_ (.Y(_1253_),
    .B(net451),
    .A_N(net1084));
 sg13g2_a21oi_1 _5603_ (.A1(_1181_),
    .A2(_1253_),
    .Y(_1254_),
    .B1(net1078));
 sg13g2_nor2b_1 _5604_ (.A(net1040),
    .B_N(net1067),
    .Y(_1255_));
 sg13g2_a21oi_1 _5605_ (.A1(net1040),
    .A2(net451),
    .Y(_1256_),
    .B1(_1255_));
 sg13g2_o21ai_1 _5606_ (.B1(net1344),
    .Y(_1257_),
    .A1(net934),
    .A2(_1256_));
 sg13g2_or2_1 _5607_ (.X(_1258_),
    .B(net506),
    .A(net1344));
 sg13g2_o21ai_1 _5608_ (.B1(_1258_),
    .Y(_1259_),
    .A1(_1254_),
    .A2(_1257_));
 sg13g2_inv_1 _5609_ (.Y(_0137_),
    .A(_1259_));
 sg13g2_mux2_1 _5610_ (.A0(\s0.data_out[9][3] ),
    .A1(\s0.data_out[10][3] ),
    .S(net1087),
    .X(_1260_));
 sg13g2_nand2_1 _5611_ (.Y(_1261_),
    .A(net934),
    .B(_1260_));
 sg13g2_and2_1 _5612_ (.A(net1036),
    .B(\s0.data_out[9][3] ),
    .X(_1262_));
 sg13g2_nor2b_1 _5613_ (.A(net1036),
    .B_N(net1062),
    .Y(_1263_));
 sg13g2_o21ai_1 _5614_ (.B1(net1079),
    .Y(_1264_),
    .A1(_1262_),
    .A2(_1263_));
 sg13g2_nand3_1 _5615_ (.B(_1261_),
    .C(_1264_),
    .A(net1341),
    .Y(_1265_));
 sg13g2_o21ai_1 _5616_ (.B1(_1265_),
    .Y(_1266_),
    .A1(net1341),
    .A2(net436));
 sg13g2_inv_1 _5617_ (.Y(_0138_),
    .A(_1266_));
 sg13g2_mux2_1 _5618_ (.A0(\s0.data_out[9][4] ),
    .A1(\s0.data_out[10][4] ),
    .S(net1086),
    .X(_1267_));
 sg13g2_nand2_1 _5619_ (.Y(_1268_),
    .A(net934),
    .B(_1267_));
 sg13g2_and2_1 _5620_ (.A(net1040),
    .B(\s0.data_out[9][4] ),
    .X(_1269_));
 sg13g2_nor2b_1 _5621_ (.A(net1040),
    .B_N(net1060),
    .Y(_1270_));
 sg13g2_o21ai_1 _5622_ (.B1(net1082),
    .Y(_1271_),
    .A1(_1269_),
    .A2(_1270_));
 sg13g2_nand3_1 _5623_ (.B(_1268_),
    .C(_1271_),
    .A(net1344),
    .Y(_1272_));
 sg13g2_o21ai_1 _5624_ (.B1(_1272_),
    .Y(_1273_),
    .A1(net1344),
    .A2(net429));
 sg13g2_inv_1 _5625_ (.Y(_0139_),
    .A(_1273_));
 sg13g2_o21ai_1 _5626_ (.B1(_1214_),
    .Y(_1274_),
    .A1(net1087),
    .A2(_2490_));
 sg13g2_nand2_1 _5627_ (.Y(_1275_),
    .A(_2454_),
    .B(_1274_));
 sg13g2_nor2_1 _5628_ (.A(net919),
    .B(_2490_),
    .Y(_1276_));
 sg13g2_nor2b_1 _5629_ (.A(net1038),
    .B_N(net1055),
    .Y(_1277_));
 sg13g2_o21ai_1 _5630_ (.B1(net1082),
    .Y(_1278_),
    .A1(_1276_),
    .A2(_1277_));
 sg13g2_nand3_1 _5631_ (.B(_1275_),
    .C(_1278_),
    .A(net1346),
    .Y(_1279_));
 sg13g2_o21ai_1 _5632_ (.B1(_1279_),
    .Y(_1280_),
    .A1(net1346),
    .A2(net481));
 sg13g2_inv_1 _5633_ (.Y(_0140_),
    .A(_1280_));
 sg13g2_nand2b_1 _5634_ (.Y(_1281_),
    .B(\s0.data_out[9][6] ),
    .A_N(net1086));
 sg13g2_a21oi_1 _5635_ (.A1(_1203_),
    .A2(_1281_),
    .Y(_1282_),
    .B1(net1082));
 sg13g2_nor2b_1 _5636_ (.A(net1039),
    .B_N(net1051),
    .Y(_1283_));
 sg13g2_a21oi_1 _5637_ (.A1(net1038),
    .A2(\s0.data_out[9][6] ),
    .Y(_1284_),
    .B1(_1283_));
 sg13g2_o21ai_1 _5638_ (.B1(net1346),
    .Y(_1285_),
    .A1(net934),
    .A2(_1284_));
 sg13g2_or2_1 _5639_ (.X(_1286_),
    .B(net521),
    .A(net1346));
 sg13g2_o21ai_1 _5640_ (.B1(_1286_),
    .Y(_1287_),
    .A1(_1282_),
    .A2(_1285_));
 sg13g2_inv_1 _5641_ (.Y(_0141_),
    .A(net522));
 sg13g2_nand2b_1 _5642_ (.Y(_1288_),
    .B(\s0.data_out[9][7] ),
    .A_N(net1086));
 sg13g2_a21oi_1 _5643_ (.A1(_1199_),
    .A2(_1288_),
    .Y(_1289_),
    .B1(net1083));
 sg13g2_nor2b_1 _5644_ (.A(net1039),
    .B_N(net1047),
    .Y(_1290_));
 sg13g2_a21oi_1 _5645_ (.A1(net1038),
    .A2(\s0.data_out[9][7] ),
    .Y(_1291_),
    .B1(_1290_));
 sg13g2_o21ai_1 _5646_ (.B1(net1347),
    .Y(_1292_),
    .A1(net934),
    .A2(_1291_));
 sg13g2_or2_1 _5647_ (.X(_1293_),
    .B(net531),
    .A(net1346));
 sg13g2_o21ai_1 _5648_ (.B1(_1293_),
    .Y(_1294_),
    .A1(_1289_),
    .A2(_1292_));
 sg13g2_inv_1 _5649_ (.Y(_0142_),
    .A(net532));
 sg13g2_mux2_1 _5650_ (.A0(\s0.data_out[10][2] ),
    .A1(\s0.data_out[9][2] ),
    .S(net1043),
    .X(_1295_));
 sg13g2_a21o_1 _5651_ (.A2(_1295_),
    .A1(net1040),
    .B1(_1255_),
    .X(_1296_));
 sg13g2_a21oi_1 _5652_ (.A1(net1079),
    .A2(_1296_),
    .Y(_1297_),
    .B1(_1254_));
 sg13g2_or2_1 _5653_ (.X(_1298_),
    .B(_1297_),
    .A(net1270));
 sg13g2_mux2_1 _5654_ (.A0(\s0.data_out[10][1] ),
    .A1(\s0.data_out[9][1] ),
    .S(net1041),
    .X(_1299_));
 sg13g2_a21oi_1 _5655_ (.A1(net1036),
    .A2(_1299_),
    .Y(_1300_),
    .B1(_1249_));
 sg13g2_nand2b_1 _5656_ (.Y(_1301_),
    .B(net1078),
    .A_N(_1300_));
 sg13g2_and2_1 _5657_ (.A(_1247_),
    .B(_1301_),
    .X(_1302_));
 sg13g2_mux2_1 _5658_ (.A0(\s0.data_out[10][0] ),
    .A1(\s0.data_out[9][0] ),
    .S(net1041),
    .X(_1303_));
 sg13g2_a21oi_1 _5659_ (.A1(net1035),
    .A2(_1303_),
    .Y(_1304_),
    .B1(_1242_));
 sg13g2_nand2b_1 _5660_ (.Y(_1305_),
    .B(net1078),
    .A_N(_1304_));
 sg13g2_a221oi_1 _5661_ (.B2(_1240_),
    .C1(net1283),
    .B1(_1305_),
    .A1(net1278),
    .Y(_1306_),
    .A2(_1302_));
 sg13g2_o21ai_1 _5662_ (.B1(_1298_),
    .Y(_1307_),
    .A1(net1278),
    .A2(_1302_));
 sg13g2_mux2_1 _5663_ (.A0(\s0.data_out[10][3] ),
    .A1(\s0.data_out[9][3] ),
    .S(net1041),
    .X(_1308_));
 sg13g2_a21oi_1 _5664_ (.A1(net1036),
    .A2(_1308_),
    .Y(_1309_),
    .B1(_1263_));
 sg13g2_nand2b_1 _5665_ (.Y(_1310_),
    .B(net1079),
    .A_N(_1309_));
 sg13g2_and2_1 _5666_ (.A(_1261_),
    .B(_1310_),
    .X(_1311_));
 sg13g2_a22oi_1 _5667_ (.Y(_1312_),
    .B1(_1311_),
    .B2(net1265),
    .A2(_1297_),
    .A1(net1270));
 sg13g2_o21ai_1 _5668_ (.B1(_1312_),
    .Y(_1313_),
    .A1(_1306_),
    .A2(_1307_));
 sg13g2_nand2_1 _5669_ (.Y(_1314_),
    .A(net1043),
    .B(net565));
 sg13g2_mux2_1 _5670_ (.A0(\s0.data_out[10][7] ),
    .A1(\s0.data_out[9][7] ),
    .S(net1043),
    .X(_1315_));
 sg13g2_a21o_1 _5671_ (.A2(_1315_),
    .A1(net1039),
    .B1(_1290_),
    .X(_1316_));
 sg13g2_a21oi_1 _5672_ (.A1(net1083),
    .A2(_1316_),
    .Y(_1317_),
    .B1(_1289_));
 sg13g2_nand2_1 _5673_ (.Y(_1318_),
    .A(net1041),
    .B(net542));
 sg13g2_mux2_1 _5674_ (.A0(\s0.data_out[10][6] ),
    .A1(\s0.data_out[9][6] ),
    .S(net1043),
    .X(_1319_));
 sg13g2_a21o_1 _5675_ (.A2(_1319_),
    .A1(net1039),
    .B1(_1283_),
    .X(_1320_));
 sg13g2_a21oi_1 _5676_ (.A1(net1083),
    .A2(_1320_),
    .Y(_1321_),
    .B1(_1282_));
 sg13g2_a22oi_1 _5677_ (.Y(_1322_),
    .B1(_1321_),
    .B2(net1243),
    .A2(_1317_),
    .A1(net1237));
 sg13g2_inv_1 _5678_ (.Y(_1323_),
    .A(_1322_));
 sg13g2_nor2_1 _5679_ (.A(net1243),
    .B(_1321_),
    .Y(_1324_));
 sg13g2_or2_1 _5680_ (.X(_1325_),
    .B(_1317_),
    .A(net1237));
 sg13g2_nand2_1 _5681_ (.Y(_1326_),
    .A(_1322_),
    .B(_1325_));
 sg13g2_nor2_1 _5682_ (.A(_1324_),
    .B(_1326_),
    .Y(_1327_));
 sg13g2_mux2_1 _5683_ (.A0(\s0.data_out[10][4] ),
    .A1(\s0.data_out[9][4] ),
    .S(net1043),
    .X(_1328_));
 sg13g2_a21oi_1 _5684_ (.A1(net1040),
    .A2(_1328_),
    .Y(_1329_),
    .B1(_1270_));
 sg13g2_nand2b_1 _5685_ (.Y(_1330_),
    .B(net1082),
    .A_N(_1329_));
 sg13g2_nand3_1 _5686_ (.B(_1268_),
    .C(_1330_),
    .A(net1257),
    .Y(_1331_));
 sg13g2_mux2_1 _5687_ (.A0(\s0.data_out[10][5] ),
    .A1(\s0.data_out[9][5] ),
    .S(net1043),
    .X(_1332_));
 sg13g2_a21oi_1 _5688_ (.A1(net1038),
    .A2(_1332_),
    .Y(_1333_),
    .B1(_1277_));
 sg13g2_nand2b_1 _5689_ (.Y(_1334_),
    .B(net1082),
    .A_N(_1333_));
 sg13g2_nand3_1 _5690_ (.B(_1275_),
    .C(_1334_),
    .A(net1252),
    .Y(_1335_));
 sg13g2_nand2_1 _5691_ (.Y(_1336_),
    .A(_1331_),
    .B(_1335_));
 sg13g2_a21oi_1 _5692_ (.A1(_1268_),
    .A2(_1330_),
    .Y(_1337_),
    .B1(net1257));
 sg13g2_nor2_1 _5693_ (.A(net1266),
    .B(_1311_),
    .Y(_1338_));
 sg13g2_a21oi_1 _5694_ (.A1(_1275_),
    .A2(_1334_),
    .Y(_1339_),
    .B1(net1251));
 sg13g2_nor4_1 _5695_ (.A(_1336_),
    .B(_1337_),
    .C(_1338_),
    .D(_1339_),
    .Y(_1340_));
 sg13g2_nand3_1 _5696_ (.B(_1327_),
    .C(_1340_),
    .A(_1313_),
    .Y(_1341_));
 sg13g2_o21ai_1 _5697_ (.B1(_1335_),
    .Y(_1342_),
    .A1(_1331_),
    .A2(_1339_));
 sg13g2_a221oi_1 _5698_ (.B2(_1342_),
    .C1(_1233_),
    .B1(_1327_),
    .A1(_1323_),
    .Y(_1343_),
    .A2(_1325_));
 sg13g2_or2_1 _5699_ (.X(_1344_),
    .B(net1210),
    .A(net315));
 sg13g2_a21oi_1 _5700_ (.A1(_1341_),
    .A2(_1343_),
    .Y(_0143_),
    .B1(_1344_));
 sg13g2_mux2_1 _5701_ (.A0(net1073),
    .A1(net1281),
    .S(net1223),
    .X(_0144_));
 sg13g2_mux2_1 _5702_ (.A0(net1069),
    .A1(net1273),
    .S(net1224),
    .X(_0145_));
 sg13g2_nor2_1 _5703_ (.A(net1224),
    .B(net1065),
    .Y(_1345_));
 sg13g2_a21oi_1 _5704_ (.A1(net1223),
    .A2(net1211),
    .Y(_0146_),
    .B1(_1345_));
 sg13g2_mux2_1 _5705_ (.A0(net1061),
    .A1(net1260),
    .S(net1224),
    .X(_0147_));
 sg13g2_nor2_1 _5706_ (.A(net1224),
    .B(net1057),
    .Y(_1346_));
 sg13g2_a21oi_1 _5707_ (.A1(net1223),
    .A2(net1214),
    .Y(_0148_),
    .B1(_1346_));
 sg13g2_mux2_1 _5708_ (.A0(net1053),
    .A1(net1246),
    .S(net1223),
    .X(_0149_));
 sg13g2_nor2_1 _5709_ (.A(net1223),
    .B(net1049),
    .Y(_1347_));
 sg13g2_a21oi_1 _5710_ (.A1(net1223),
    .A2(_2474_),
    .Y(_0150_),
    .B1(_1347_));
 sg13g2_mux2_1 _5711_ (.A0(net1045),
    .A1(net1231),
    .S(net1223),
    .X(_0151_));
 sg13g2_o21ai_1 _5712_ (.B1(net1037),
    .Y(_1348_),
    .A1(net1230),
    .A2(net1028));
 sg13g2_nor2b_1 _5713_ (.A(net1230),
    .B_N(net1033),
    .Y(_1349_));
 sg13g2_nor2_1 _5714_ (.A(_1348_),
    .B(_1349_),
    .Y(_1350_));
 sg13g2_inv_1 _5715_ (.Y(_1351_),
    .A(_1350_));
 sg13g2_o21ai_1 _5716_ (.B1(_1351_),
    .Y(_1352_),
    .A1(net1038),
    .A2(_1230_));
 sg13g2_or2_1 _5717_ (.X(_1353_),
    .B(net1033),
    .A(net398));
 sg13g2_o21ai_1 _5718_ (.B1(net920),
    .Y(_1354_),
    .A1(net398),
    .A2(net1042));
 sg13g2_o21ai_1 _5719_ (.B1(_1354_),
    .Y(_1355_),
    .A1(net1028),
    .A2(_1348_));
 sg13g2_a21oi_1 _5720_ (.A1(_1350_),
    .A2(_1353_),
    .Y(_1356_),
    .B1(_1355_));
 sg13g2_o21ai_1 _5721_ (.B1(net1346),
    .Y(_1357_),
    .A1(net453),
    .A2(_1352_));
 sg13g2_nor2_1 _5722_ (.A(_1356_),
    .B(_1357_),
    .Y(_0152_));
 sg13g2_nor2_1 _5723_ (.A(net1221),
    .B(_1352_),
    .Y(_0153_));
 sg13g2_mux2_1 _5724_ (.A0(\s0.data_out[8][0] ),
    .A1(\s0.data_out[9][0] ),
    .S(net1041),
    .X(_1358_));
 sg13g2_nand2_1 _5725_ (.Y(_1359_),
    .A(net919),
    .B(_1358_));
 sg13g2_and2_1 _5726_ (.A(net1023),
    .B(\s0.data_out[8][0] ),
    .X(_1360_));
 sg13g2_nor2b_1 _5727_ (.A(net1024),
    .B_N(net1075),
    .Y(_1361_));
 sg13g2_o21ai_1 _5728_ (.B1(net1035),
    .Y(_1362_),
    .A1(_1360_),
    .A2(_1361_));
 sg13g2_nand3_1 _5729_ (.B(_1359_),
    .C(_1362_),
    .A(net1340),
    .Y(_1363_));
 sg13g2_o21ai_1 _5730_ (.B1(_1363_),
    .Y(_1364_),
    .A1(net1340),
    .A2(net428));
 sg13g2_inv_1 _5731_ (.Y(_0154_),
    .A(_1364_));
 sg13g2_mux2_1 _5732_ (.A0(\s0.data_out[8][1] ),
    .A1(\s0.data_out[9][1] ),
    .S(net1041),
    .X(_1365_));
 sg13g2_nand2_1 _5733_ (.Y(_1366_),
    .A(net919),
    .B(_1365_));
 sg13g2_and2_1 _5734_ (.A(net1030),
    .B(\s0.data_out[8][1] ),
    .X(_1367_));
 sg13g2_nor2b_1 _5735_ (.A(net1030),
    .B_N(net1071),
    .Y(_1368_));
 sg13g2_o21ai_1 _5736_ (.B1(net1035),
    .Y(_1369_),
    .A1(_1367_),
    .A2(_1368_));
 sg13g2_nand3_1 _5737_ (.B(_1366_),
    .C(_1369_),
    .A(net1341),
    .Y(_1370_));
 sg13g2_o21ai_1 _5738_ (.B1(_1370_),
    .Y(_1371_),
    .A1(net1340),
    .A2(net405));
 sg13g2_inv_1 _5739_ (.Y(_0155_),
    .A(_1371_));
 sg13g2_mux2_1 _5740_ (.A0(\s0.data_out[8][2] ),
    .A1(\s0.data_out[9][2] ),
    .S(net1041),
    .X(_1372_));
 sg13g2_nand2_1 _5741_ (.Y(_1373_),
    .A(net919),
    .B(_1372_));
 sg13g2_and2_1 _5742_ (.A(net1024),
    .B(net608),
    .X(_1374_));
 sg13g2_nor2b_1 _5743_ (.A(net1030),
    .B_N(net1067),
    .Y(_1375_));
 sg13g2_o21ai_1 _5744_ (.B1(net1036),
    .Y(_1376_),
    .A1(_1374_),
    .A2(_1375_));
 sg13g2_nand3_1 _5745_ (.B(_1373_),
    .C(_1376_),
    .A(net1340),
    .Y(_1377_));
 sg13g2_o21ai_1 _5746_ (.B1(net609),
    .Y(_1378_),
    .A1(net1340),
    .A2(net451));
 sg13g2_inv_1 _5747_ (.Y(_0156_),
    .A(_1378_));
 sg13g2_mux2_1 _5748_ (.A0(\s0.data_out[8][3] ),
    .A1(\s0.data_out[9][3] ),
    .S(net1041),
    .X(_1379_));
 sg13g2_nand2_1 _5749_ (.Y(_1380_),
    .A(net919),
    .B(_1379_));
 sg13g2_and2_1 _5750_ (.A(net1030),
    .B(\s0.data_out[8][3] ),
    .X(_1381_));
 sg13g2_nor2b_1 _5751_ (.A(net1030),
    .B_N(net1063),
    .Y(_1382_));
 sg13g2_o21ai_1 _5752_ (.B1(net1035),
    .Y(_1383_),
    .A1(_1381_),
    .A2(_1382_));
 sg13g2_nand3_1 _5753_ (.B(_1380_),
    .C(_1383_),
    .A(net1341),
    .Y(_1384_));
 sg13g2_o21ai_1 _5754_ (.B1(_1384_),
    .Y(_1385_),
    .A1(net1340),
    .A2(net400));
 sg13g2_inv_1 _5755_ (.Y(_0157_),
    .A(_1385_));
 sg13g2_mux2_1 _5756_ (.A0(\s0.data_out[8][4] ),
    .A1(\s0.data_out[9][4] ),
    .S(net1042),
    .X(_1386_));
 sg13g2_nand2_1 _5757_ (.Y(_1387_),
    .A(net919),
    .B(_1386_));
 sg13g2_and2_1 _5758_ (.A(net1027),
    .B(\s0.data_out[8][4] ),
    .X(_1388_));
 sg13g2_nor2b_1 _5759_ (.A(net1027),
    .B_N(net1059),
    .Y(_1389_));
 sg13g2_o21ai_1 _5760_ (.B1(net1037),
    .Y(_1390_),
    .A1(_1388_),
    .A2(_1389_));
 sg13g2_nand3_1 _5761_ (.B(_1387_),
    .C(_1390_),
    .A(net1343),
    .Y(_1391_));
 sg13g2_o21ai_1 _5762_ (.B1(_1391_),
    .Y(_1392_),
    .A1(net1342),
    .A2(net442));
 sg13g2_inv_1 _5763_ (.Y(_0158_),
    .A(_1392_));
 sg13g2_mux2_1 _5764_ (.A0(\s0.data_out[8][5] ),
    .A1(\s0.data_out[9][5] ),
    .S(net1042),
    .X(_1393_));
 sg13g2_nand2_1 _5765_ (.Y(_1394_),
    .A(net920),
    .B(_1393_));
 sg13g2_and2_1 _5766_ (.A(net1029),
    .B(net610),
    .X(_1395_));
 sg13g2_nor2b_1 _5767_ (.A(net1027),
    .B_N(net1055),
    .Y(_1396_));
 sg13g2_o21ai_1 _5768_ (.B1(net1037),
    .Y(_1397_),
    .A1(_1395_),
    .A2(_1396_));
 sg13g2_nand3_1 _5769_ (.B(_1394_),
    .C(_1397_),
    .A(net1342),
    .Y(_1398_));
 sg13g2_o21ai_1 _5770_ (.B1(_1398_),
    .Y(_1399_),
    .A1(net1343),
    .A2(net385));
 sg13g2_inv_1 _5771_ (.Y(_0159_),
    .A(_1399_));
 sg13g2_nand2b_1 _5772_ (.Y(_1400_),
    .B(\s0.data_out[8][6] ),
    .A_N(net1042));
 sg13g2_a21oi_1 _5773_ (.A1(_1318_),
    .A2(_1400_),
    .Y(_1401_),
    .B1(net1037));
 sg13g2_nor2b_1 _5774_ (.A(net1027),
    .B_N(net1052),
    .Y(_1402_));
 sg13g2_a21oi_1 _5775_ (.A1(net1027),
    .A2(\s0.data_out[8][6] ),
    .Y(_1403_),
    .B1(_1402_));
 sg13g2_o21ai_1 _5776_ (.B1(net1343),
    .Y(_1404_),
    .A1(net920),
    .A2(_1403_));
 sg13g2_or2_1 _5777_ (.X(_1405_),
    .B(net542),
    .A(net1342));
 sg13g2_o21ai_1 _5778_ (.B1(_1405_),
    .Y(_1406_),
    .A1(_1401_),
    .A2(_1404_));
 sg13g2_inv_1 _5779_ (.Y(_0160_),
    .A(net543));
 sg13g2_nand2b_1 _5780_ (.Y(_1407_),
    .B(\s0.data_out[8][7] ),
    .A_N(net1043));
 sg13g2_a21oi_1 _5781_ (.A1(_1314_),
    .A2(_1407_),
    .Y(_1408_),
    .B1(net1038));
 sg13g2_nor2b_1 _5782_ (.A(net1027),
    .B_N(net1047),
    .Y(_1409_));
 sg13g2_a21oi_1 _5783_ (.A1(net1028),
    .A2(\s0.data_out[8][7] ),
    .Y(_1410_),
    .B1(_1409_));
 sg13g2_o21ai_1 _5784_ (.B1(net1343),
    .Y(_1411_),
    .A1(net920),
    .A2(_1410_));
 sg13g2_or2_1 _5785_ (.X(_1412_),
    .B(net565),
    .A(net1346));
 sg13g2_o21ai_1 _5786_ (.B1(_1412_),
    .Y(_1413_),
    .A1(_1408_),
    .A2(_1411_));
 sg13g2_inv_1 _5787_ (.Y(_0161_),
    .A(net566));
 sg13g2_nand2_1 _5788_ (.Y(_1414_),
    .A(net1031),
    .B(net487));
 sg13g2_o21ai_1 _5789_ (.B1(_1414_),
    .Y(_1415_),
    .A1(net1031),
    .A2(_2489_));
 sg13g2_a21oi_1 _5790_ (.A1(net1030),
    .A2(_1415_),
    .Y(_1416_),
    .B1(_1375_));
 sg13g2_o21ai_1 _5791_ (.B1(_1373_),
    .Y(_1417_),
    .A1(net919),
    .A2(_1416_));
 sg13g2_nand2_1 _5792_ (.Y(_1418_),
    .A(net1031),
    .B(net526));
 sg13g2_mux2_1 _5793_ (.A0(\s0.data_out[9][1] ),
    .A1(\s0.data_out[8][1] ),
    .S(net1034),
    .X(_1419_));
 sg13g2_a21oi_1 _5794_ (.A1(net1030),
    .A2(_1419_),
    .Y(_1420_),
    .B1(_1368_));
 sg13g2_nand2b_1 _5795_ (.Y(_1421_),
    .B(net1035),
    .A_N(_1420_));
 sg13g2_nand3_1 _5796_ (.B(_1366_),
    .C(_1421_),
    .A(net1280),
    .Y(_1422_));
 sg13g2_mux2_1 _5797_ (.A0(\s0.data_out[9][0] ),
    .A1(\s0.data_out[8][0] ),
    .S(net1031),
    .X(_1423_));
 sg13g2_a21oi_1 _5798_ (.A1(net1024),
    .A2(_1423_),
    .Y(_1424_),
    .B1(_1361_));
 sg13g2_o21ai_1 _5799_ (.B1(_1359_),
    .Y(_1425_),
    .A1(net919),
    .A2(_1424_));
 sg13g2_nor2b_1 _5800_ (.A(net1283),
    .B_N(_1425_),
    .Y(_1426_));
 sg13g2_a21oi_1 _5801_ (.A1(_1366_),
    .A2(_1421_),
    .Y(_1427_),
    .B1(net1279));
 sg13g2_a221oi_1 _5802_ (.B2(_1426_),
    .C1(_1427_),
    .B1(_1422_),
    .A1(net1213),
    .Y(_1428_),
    .A2(_1417_));
 sg13g2_mux2_1 _5803_ (.A0(\s0.data_out[9][3] ),
    .A1(\s0.data_out[8][3] ),
    .S(net1034),
    .X(_1429_));
 sg13g2_a21oi_1 _5804_ (.A1(net1030),
    .A2(_1429_),
    .Y(_1430_),
    .B1(_1382_));
 sg13g2_nand2b_1 _5805_ (.Y(_1431_),
    .B(net1035),
    .A_N(_1430_));
 sg13g2_and2_1 _5806_ (.A(_1380_),
    .B(_1431_),
    .X(_1432_));
 sg13g2_nand2_1 _5807_ (.Y(_1433_),
    .A(net1266),
    .B(_1432_));
 sg13g2_or2_1 _5808_ (.X(_1434_),
    .B(_1417_),
    .A(net1213));
 sg13g2_nand3b_1 _5809_ (.B(_1433_),
    .C(_1434_),
    .Y(_1435_),
    .A_N(_1428_));
 sg13g2_nand2_1 _5810_ (.Y(_1436_),
    .A(net1032),
    .B(net595));
 sg13g2_mux2_1 _5811_ (.A0(\s0.data_out[9][7] ),
    .A1(\s0.data_out[8][7] ),
    .S(net1032),
    .X(_1437_));
 sg13g2_a21o_1 _5812_ (.A2(_1437_),
    .A1(net1028),
    .B1(_1409_),
    .X(_1438_));
 sg13g2_a21oi_1 _5813_ (.A1(net1038),
    .A2(_1438_),
    .Y(_1439_),
    .B1(_1408_));
 sg13g2_nand2_1 _5814_ (.Y(_1440_),
    .A(net1032),
    .B(net587));
 sg13g2_mux2_1 _5815_ (.A0(\s0.data_out[9][6] ),
    .A1(\s0.data_out[8][6] ),
    .S(net1033),
    .X(_1441_));
 sg13g2_a21o_1 _5816_ (.A2(_1441_),
    .A1(net1028),
    .B1(_1402_),
    .X(_1442_));
 sg13g2_a21oi_1 _5817_ (.A1(net1037),
    .A2(_1442_),
    .Y(_1443_),
    .B1(_1401_));
 sg13g2_a22oi_1 _5818_ (.Y(_1444_),
    .B1(_1443_),
    .B2(net1243),
    .A2(_1439_),
    .A1(net1237));
 sg13g2_inv_1 _5819_ (.Y(_1445_),
    .A(_1444_));
 sg13g2_nor2_1 _5820_ (.A(net1243),
    .B(_1443_),
    .Y(_1446_));
 sg13g2_or2_1 _5821_ (.X(_1447_),
    .B(_1439_),
    .A(net1237));
 sg13g2_nand2_1 _5822_ (.Y(_1448_),
    .A(_1444_),
    .B(_1447_));
 sg13g2_nor2_1 _5823_ (.A(_1446_),
    .B(_1448_),
    .Y(_1449_));
 sg13g2_nand2_1 _5824_ (.Y(_1450_),
    .A(net1033),
    .B(net482));
 sg13g2_o21ai_1 _5825_ (.B1(_1450_),
    .Y(_1451_),
    .A1(net1033),
    .A2(_2490_));
 sg13g2_a21oi_1 _5826_ (.A1(net1027),
    .A2(_1451_),
    .Y(_1452_),
    .B1(_1396_));
 sg13g2_nand2b_1 _5827_ (.Y(_1453_),
    .B(net1037),
    .A_N(_1452_));
 sg13g2_nand3_1 _5828_ (.B(_1394_),
    .C(_1453_),
    .A(net1252),
    .Y(_1454_));
 sg13g2_mux2_1 _5829_ (.A0(\s0.data_out[9][4] ),
    .A1(\s0.data_out[8][4] ),
    .S(net1033),
    .X(_1455_));
 sg13g2_a21oi_1 _5830_ (.A1(net1027),
    .A2(_1455_),
    .Y(_1456_),
    .B1(_1389_));
 sg13g2_nand2b_1 _5831_ (.Y(_1457_),
    .B(net343),
    .A_N(_1456_));
 sg13g2_nand3_1 _5832_ (.B(_1387_),
    .C(_1457_),
    .A(net1257),
    .Y(_1458_));
 sg13g2_and2_1 _5833_ (.A(_1454_),
    .B(_1458_),
    .X(_1459_));
 sg13g2_a21oi_1 _5834_ (.A1(_1394_),
    .A2(_1453_),
    .Y(_1460_),
    .B1(net1252));
 sg13g2_nor2_1 _5835_ (.A(net1266),
    .B(_1432_),
    .Y(_1461_));
 sg13g2_a21oi_1 _5836_ (.A1(_1387_),
    .A2(_1457_),
    .Y(_1462_),
    .B1(net1257));
 sg13g2_nor3_1 _5837_ (.A(_1460_),
    .B(_1461_),
    .C(_1462_),
    .Y(_1463_));
 sg13g2_nand4_1 _5838_ (.B(_1449_),
    .C(_1459_),
    .A(_1435_),
    .Y(_1464_),
    .D(_1463_));
 sg13g2_o21ai_1 _5839_ (.B1(_1454_),
    .Y(_1465_),
    .A1(_1458_),
    .A2(_1460_));
 sg13g2_a221oi_1 _5840_ (.B2(_1465_),
    .C1(_1352_),
    .B1(_1449_),
    .A1(_1445_),
    .Y(_1466_),
    .A2(_1447_));
 sg13g2_or2_1 _5841_ (.X(_1467_),
    .B(net1210),
    .A(net314));
 sg13g2_a21oi_1 _5842_ (.A1(_1464_),
    .A2(_1466_),
    .Y(_0162_),
    .B1(_1467_));
 sg13g2_and2_1 _5843_ (.A(net1329),
    .B(net307),
    .X(_0163_));
 sg13g2_o21ai_1 _5844_ (.B1(net1025),
    .Y(_1468_),
    .A1(net1230),
    .A2(net1016));
 sg13g2_a21oi_1 _5845_ (.A1(_2449_),
    .A2(net1021),
    .Y(_1469_),
    .B1(_1468_));
 sg13g2_inv_1 _5846_ (.Y(_1470_),
    .A(_1469_));
 sg13g2_o21ai_1 _5847_ (.B1(_1470_),
    .Y(_1471_),
    .A1(net1029),
    .A2(_1349_));
 sg13g2_o21ai_1 _5848_ (.B1(_1469_),
    .Y(_1472_),
    .A1(net326),
    .A2(net1021));
 sg13g2_nor2_1 _5849_ (.A(net1016),
    .B(_1468_),
    .Y(_1473_));
 sg13g2_o21ai_1 _5850_ (.B1(net918),
    .Y(_1474_),
    .A1(net326),
    .A2(net1032));
 sg13g2_nor2b_1 _5851_ (.A(_1473_),
    .B_N(_1474_),
    .Y(_1475_));
 sg13g2_o21ai_1 _5852_ (.B1(net1342),
    .Y(_1476_),
    .A1(net398),
    .A2(_1471_));
 sg13g2_a21oi_1 _5853_ (.A1(_1472_),
    .A2(_1475_),
    .Y(_0164_),
    .B1(_1476_));
 sg13g2_nor2_1 _5854_ (.A(net1221),
    .B(_1471_),
    .Y(_0165_));
 sg13g2_mux2_1 _5855_ (.A0(\s0.data_out[7][0] ),
    .A1(\s0.data_out[8][0] ),
    .S(net1031),
    .X(_1477_));
 sg13g2_nand2_1 _5856_ (.Y(_1478_),
    .A(net918),
    .B(_1477_));
 sg13g2_and2_1 _5857_ (.A(net1012),
    .B(\s0.data_out[7][0] ),
    .X(_1479_));
 sg13g2_nor2b_1 _5858_ (.A(net1013),
    .B_N(net1075),
    .Y(_1480_));
 sg13g2_o21ai_1 _5859_ (.B1(net1023),
    .Y(_1481_),
    .A1(_1479_),
    .A2(_1480_));
 sg13g2_nand3_1 _5860_ (.B(_1478_),
    .C(_1481_),
    .A(net1328),
    .Y(_1482_));
 sg13g2_o21ai_1 _5861_ (.B1(_1482_),
    .Y(_1483_),
    .A1(net1328),
    .A2(net390));
 sg13g2_inv_1 _5862_ (.Y(_0166_),
    .A(_1483_));
 sg13g2_nand2b_1 _5863_ (.Y(_1484_),
    .B(net419),
    .A_N(net1031));
 sg13g2_a21oi_1 _5864_ (.A1(_1418_),
    .A2(_1484_),
    .Y(_1485_),
    .B1(net1023));
 sg13g2_nor2b_1 _5865_ (.A(net1013),
    .B_N(net1071),
    .Y(_1486_));
 sg13g2_a21oi_1 _5866_ (.A1(net1013),
    .A2(net419),
    .Y(_1487_),
    .B1(_1486_));
 sg13g2_o21ai_1 _5867_ (.B1(net1328),
    .Y(_1488_),
    .A1(net918),
    .A2(_1487_));
 sg13g2_or2_1 _5868_ (.X(_1489_),
    .B(net526),
    .A(net1328));
 sg13g2_o21ai_1 _5869_ (.B1(_1489_),
    .Y(_1490_),
    .A1(_1485_),
    .A2(_1488_));
 sg13g2_inv_1 _5870_ (.Y(_0167_),
    .A(_1490_));
 sg13g2_nand2b_1 _5871_ (.Y(_1491_),
    .B(net467),
    .A_N(net1031));
 sg13g2_a21oi_1 _5872_ (.A1(_1414_),
    .A2(_1491_),
    .Y(_1492_),
    .B1(net1024));
 sg13g2_nor2b_1 _5873_ (.A(net1013),
    .B_N(net1067),
    .Y(_1493_));
 sg13g2_a21oi_1 _5874_ (.A1(net1013),
    .A2(net467),
    .Y(_1494_),
    .B1(_1493_));
 sg13g2_o21ai_1 _5875_ (.B1(net1328),
    .Y(_1495_),
    .A1(net918),
    .A2(_1494_));
 sg13g2_or2_1 _5876_ (.X(_1496_),
    .B(net487),
    .A(net1328));
 sg13g2_o21ai_1 _5877_ (.B1(_1496_),
    .Y(_1497_),
    .A1(_1492_),
    .A2(_1495_));
 sg13g2_inv_1 _5878_ (.Y(_0168_),
    .A(_1497_));
 sg13g2_mux2_1 _5879_ (.A0(\s0.data_out[7][3] ),
    .A1(\s0.data_out[8][3] ),
    .S(net1031),
    .X(_1498_));
 sg13g2_nand2_1 _5880_ (.Y(_1499_),
    .A(net918),
    .B(_1498_));
 sg13g2_and2_1 _5881_ (.A(net1012),
    .B(\s0.data_out[7][3] ),
    .X(_1500_));
 sg13g2_nor2b_1 _5882_ (.A(net1014),
    .B_N(net1063),
    .Y(_1501_));
 sg13g2_o21ai_1 _5883_ (.B1(net1023),
    .Y(_1502_),
    .A1(_1500_),
    .A2(_1501_));
 sg13g2_nand3_1 _5884_ (.B(_1499_),
    .C(_1502_),
    .A(net1328),
    .Y(_1503_));
 sg13g2_o21ai_1 _5885_ (.B1(_1503_),
    .Y(_1504_),
    .A1(net1327),
    .A2(net434));
 sg13g2_inv_1 _5886_ (.Y(_0169_),
    .A(_1504_));
 sg13g2_mux2_1 _5887_ (.A0(\s0.data_out[7][4] ),
    .A1(\s0.data_out[8][4] ),
    .S(net1032),
    .X(_1505_));
 sg13g2_nand2_1 _5888_ (.Y(_1506_),
    .A(_2467_),
    .B(_1505_));
 sg13g2_and2_1 _5889_ (.A(net1016),
    .B(\s0.data_out[7][4] ),
    .X(_1507_));
 sg13g2_nor2b_1 _5890_ (.A(net1016),
    .B_N(net1059),
    .Y(_1508_));
 sg13g2_o21ai_1 _5891_ (.B1(net1025),
    .Y(_1509_),
    .A1(_1507_),
    .A2(_1508_));
 sg13g2_nand3_1 _5892_ (.B(_1506_),
    .C(_1509_),
    .A(net1330),
    .Y(_1510_));
 sg13g2_o21ai_1 _5893_ (.B1(_1510_),
    .Y(_1511_),
    .A1(net1330),
    .A2(net350));
 sg13g2_inv_1 _5894_ (.Y(_0170_),
    .A(_1511_));
 sg13g2_nand2b_1 _5895_ (.Y(_1512_),
    .B(\s0.data_out[7][5] ),
    .A_N(net1032));
 sg13g2_a21oi_1 _5896_ (.A1(_1450_),
    .A2(_1512_),
    .Y(_1513_),
    .B1(net1025));
 sg13g2_nor2b_1 _5897_ (.A(net1016),
    .B_N(net1056),
    .Y(_1514_));
 sg13g2_a21oi_1 _5898_ (.A1(net1016),
    .A2(\s0.data_out[7][5] ),
    .Y(_1515_),
    .B1(_1514_));
 sg13g2_o21ai_1 _5899_ (.B1(net1342),
    .Y(_1516_),
    .A1(net918),
    .A2(_1515_));
 sg13g2_or2_1 _5900_ (.X(_1517_),
    .B(net482),
    .A(net1342));
 sg13g2_o21ai_1 _5901_ (.B1(_1517_),
    .Y(_1518_),
    .A1(_1513_),
    .A2(_1516_));
 sg13g2_inv_1 _5902_ (.Y(_0171_),
    .A(net483));
 sg13g2_nand2b_1 _5903_ (.Y(_1519_),
    .B(net544),
    .A_N(net1032));
 sg13g2_a21oi_1 _5904_ (.A1(_1440_),
    .A2(_1519_),
    .Y(_1520_),
    .B1(net1025));
 sg13g2_nor2b_1 _5905_ (.A(net1017),
    .B_N(net1051),
    .Y(_1521_));
 sg13g2_a21oi_1 _5906_ (.A1(net1017),
    .A2(net544),
    .Y(_1522_),
    .B1(_1521_));
 sg13g2_o21ai_1 _5907_ (.B1(net1330),
    .Y(_1523_),
    .A1(net918),
    .A2(_1522_));
 sg13g2_or2_1 _5908_ (.X(_1524_),
    .B(net587),
    .A(net1330));
 sg13g2_o21ai_1 _5909_ (.B1(_1524_),
    .Y(_1525_),
    .A1(_1520_),
    .A2(_1523_));
 sg13g2_inv_1 _5910_ (.Y(_0172_),
    .A(_1525_));
 sg13g2_nand2b_1 _5911_ (.Y(_1526_),
    .B(net517),
    .A_N(net1032));
 sg13g2_a21oi_1 _5912_ (.A1(_1436_),
    .A2(_1526_),
    .Y(_1527_),
    .B1(net1026));
 sg13g2_nor2b_1 _5913_ (.A(net1017),
    .B_N(net1048),
    .Y(_1528_));
 sg13g2_a21oi_1 _5914_ (.A1(net1017),
    .A2(net517),
    .Y(_1529_),
    .B1(_1528_));
 sg13g2_o21ai_1 _5915_ (.B1(net1330),
    .Y(_1530_),
    .A1(net918),
    .A2(_1529_));
 sg13g2_or2_1 _5916_ (.X(_1531_),
    .B(net595),
    .A(net1342));
 sg13g2_o21ai_1 _5917_ (.B1(_1531_),
    .Y(_1532_),
    .A1(_1527_),
    .A2(_1530_));
 sg13g2_inv_1 _5918_ (.Y(_0173_),
    .A(net596));
 sg13g2_mux2_1 _5919_ (.A0(\s0.data_out[8][2] ),
    .A1(\s0.data_out[7][2] ),
    .S(net1019),
    .X(_1533_));
 sg13g2_a21o_1 _5920_ (.A2(_1533_),
    .A1(net1013),
    .B1(_1493_),
    .X(_1534_));
 sg13g2_a21oi_1 _5921_ (.A1(net1023),
    .A2(_1534_),
    .Y(_1535_),
    .B1(_1492_));
 sg13g2_or2_1 _5922_ (.X(_1536_),
    .B(_1535_),
    .A(net1272));
 sg13g2_mux2_1 _5923_ (.A0(\s0.data_out[8][1] ),
    .A1(\s0.data_out[7][1] ),
    .S(net1022),
    .X(_1537_));
 sg13g2_a21o_1 _5924_ (.A2(_1537_),
    .A1(net1013),
    .B1(_1486_),
    .X(_1538_));
 sg13g2_a21oi_1 _5925_ (.A1(net1023),
    .A2(_1538_),
    .Y(_1539_),
    .B1(_1485_));
 sg13g2_mux2_1 _5926_ (.A0(\s0.data_out[8][0] ),
    .A1(\s0.data_out[7][0] ),
    .S(net1019),
    .X(_1540_));
 sg13g2_a21oi_1 _5927_ (.A1(net1013),
    .A2(_1540_),
    .Y(_1541_),
    .B1(_1480_));
 sg13g2_nand2b_1 _5928_ (.Y(_1542_),
    .B(net1023),
    .A_N(_1541_));
 sg13g2_a221oi_1 _5929_ (.B2(_1478_),
    .C1(net1283),
    .B1(_1542_),
    .A1(net1278),
    .Y(_1543_),
    .A2(_1539_));
 sg13g2_o21ai_1 _5930_ (.B1(_1536_),
    .Y(_1544_),
    .A1(net1278),
    .A2(_1539_));
 sg13g2_nand2_1 _5931_ (.Y(_1545_),
    .A(net1019),
    .B(net503));
 sg13g2_mux2_1 _5932_ (.A0(\s0.data_out[8][3] ),
    .A1(\s0.data_out[7][3] ),
    .S(net1022),
    .X(_1546_));
 sg13g2_a21oi_1 _5933_ (.A1(net1014),
    .A2(_1546_),
    .Y(_1547_),
    .B1(_1501_));
 sg13g2_nand2b_1 _5934_ (.Y(_1548_),
    .B(net1023),
    .A_N(_1547_));
 sg13g2_and2_1 _5935_ (.A(_1499_),
    .B(_1548_),
    .X(_1549_));
 sg13g2_a22oi_1 _5936_ (.Y(_1550_),
    .B1(_1549_),
    .B2(net1266),
    .A2(_1535_),
    .A1(net1271));
 sg13g2_o21ai_1 _5937_ (.B1(_1550_),
    .Y(_1551_),
    .A1(_1543_),
    .A2(_1544_));
 sg13g2_nand2_1 _5938_ (.Y(_1552_),
    .A(net1020),
    .B(net517));
 sg13g2_mux2_1 _5939_ (.A0(\s0.data_out[8][7] ),
    .A1(\s0.data_out[7][7] ),
    .S(net1021),
    .X(_1553_));
 sg13g2_a21o_1 _5940_ (.A2(_1553_),
    .A1(net1017),
    .B1(_1528_),
    .X(_1554_));
 sg13g2_a21oi_1 _5941_ (.A1(net1025),
    .A2(_1554_),
    .Y(_1555_),
    .B1(_1527_));
 sg13g2_nand2_1 _5942_ (.Y(_1556_),
    .A(net1020),
    .B(net544));
 sg13g2_mux2_1 _5943_ (.A0(\s0.data_out[8][6] ),
    .A1(\s0.data_out[7][6] ),
    .S(net1021),
    .X(_1557_));
 sg13g2_a21o_1 _5944_ (.A2(_1557_),
    .A1(net1017),
    .B1(_1521_),
    .X(_1558_));
 sg13g2_a21oi_1 _5945_ (.A1(net1025),
    .A2(_1558_),
    .Y(_1559_),
    .B1(_1520_));
 sg13g2_a22oi_1 _5946_ (.Y(_1560_),
    .B1(_1559_),
    .B2(net1243),
    .A2(_1555_),
    .A1(net1237));
 sg13g2_nor2_1 _5947_ (.A(net1242),
    .B(_1559_),
    .Y(_1561_));
 sg13g2_or2_1 _5948_ (.X(_1562_),
    .B(_1555_),
    .A(net1237));
 sg13g2_nand3b_1 _5949_ (.B(_1562_),
    .C(_1560_),
    .Y(_1563_),
    .A_N(_1561_));
 sg13g2_dfrbpq_1 _5950_ (.RESET_B(net221),
    .D(_0000_),
    .Q(\s0.module0.bubble ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _5951_ (.RESET_B(net67),
    .D(net373),
    .Q(\s0.was_valid_out[21] [0]),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _5952_ (.RESET_B(net65),
    .D(_0002_),
    .Q(\s0.valid_out[21] [0]),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _5953_ (.RESET_B(net64),
    .D(net369),
    .Q(\s0.data_out[21][0] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _5954_ (.RESET_B(net63),
    .D(_0004_),
    .Q(\s0.data_out[21][1] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _5955_ (.RESET_B(net62),
    .D(_0005_),
    .Q(\s0.data_out[21][2] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _5956_ (.RESET_B(net61),
    .D(net367),
    .Q(\s0.data_out[21][3] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _5957_ (.RESET_B(net60),
    .D(net360),
    .Q(\s0.data_out[21][4] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _5958_ (.RESET_B(net59),
    .D(net362),
    .Q(\s0.data_out[21][5] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _5959_ (.RESET_B(net58),
    .D(net357),
    .Q(\s0.data_out[21][6] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _5960_ (.RESET_B(net57),
    .D(net365),
    .Q(\s0.data_out[21][7] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _5961_ (.RESET_B(net56),
    .D(_0011_),
    .Q(\s0.shift_out[21] [0]),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _5962_ (.RESET_B(net55),
    .D(_0012_),
    .Q(\s0.genblk1[20].modules.bubble ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _5963_ (.RESET_B(net54),
    .D(_0013_),
    .Q(\s0.was_valid_out[20] [0]),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _5964_ (.RESET_B(net52),
    .D(_0014_),
    .Q(\s0.valid_out[20] [0]),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _5965_ (.RESET_B(net51),
    .D(_0015_),
    .Q(\s0.data_out[20][0] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _5966_ (.RESET_B(net50),
    .D(_0016_),
    .Q(\s0.data_out[20][1] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _5967_ (.RESET_B(net49),
    .D(_0017_),
    .Q(\s0.data_out[20][2] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _5968_ (.RESET_B(net48),
    .D(_0018_),
    .Q(\s0.data_out[20][3] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _5969_ (.RESET_B(net47),
    .D(_0019_),
    .Q(\s0.data_out[20][4] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _5970_ (.RESET_B(net46),
    .D(_0020_),
    .Q(\s0.data_out[20][5] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _5971_ (.RESET_B(net45),
    .D(_0021_),
    .Q(\s0.data_out[20][6] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _5972_ (.RESET_B(net44),
    .D(_0022_),
    .Q(\s0.data_out[20][7] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _5973_ (.RESET_B(net43),
    .D(_0023_),
    .Q(\s0.shift_out[20] [0]),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _5974_ (.RESET_B(net42),
    .D(_0024_),
    .Q(\s0.genblk1[1].modules.bubble ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _5975_ (.RESET_B(net41),
    .D(net324),
    .Q(\s0.was_valid_out[19] [0]),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _5976_ (.RESET_B(net39),
    .D(_0026_),
    .Q(\s0.valid_out[19] [0]),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _5977_ (.RESET_B(net38),
    .D(_0027_),
    .Q(\s0.data_out[19][0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _5978_ (.RESET_B(net37),
    .D(_0028_),
    .Q(\s0.data_out[19][1] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _5979_ (.RESET_B(net36),
    .D(_0029_),
    .Q(\s0.data_out[19][2] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _5980_ (.RESET_B(net35),
    .D(_0030_),
    .Q(\s0.data_out[19][3] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _5981_ (.RESET_B(net34),
    .D(_0031_),
    .Q(\s0.data_out[19][4] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _5982_ (.RESET_B(net33),
    .D(_0032_),
    .Q(\s0.data_out[19][5] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _5983_ (.RESET_B(net32),
    .D(_0033_),
    .Q(\s0.data_out[19][6] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _5984_ (.RESET_B(net31),
    .D(_0034_),
    .Q(\s0.data_out[19][7] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _5985_ (.RESET_B(net30),
    .D(_0035_),
    .Q(\s0.shift_out[19] [0]),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _5986_ (.RESET_B(net29),
    .D(_0036_),
    .Q(\s0.genblk1[18].modules.bubble ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _5987_ (.RESET_B(net28),
    .D(net407),
    .Q(\s0.was_valid_out[18] [0]),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _5988_ (.RESET_B(net26),
    .D(_0038_),
    .Q(\s0.valid_out[18] [0]),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _5989_ (.RESET_B(net25),
    .D(_0039_),
    .Q(\s0.data_out[18][0] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _5990_ (.RESET_B(net24),
    .D(_0040_),
    .Q(\s0.data_out[18][1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _5991_ (.RESET_B(net23),
    .D(_0041_),
    .Q(\s0.data_out[18][2] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _5992_ (.RESET_B(net294),
    .D(_0042_),
    .Q(\s0.data_out[18][3] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _5993_ (.RESET_B(net293),
    .D(_0043_),
    .Q(\s0.data_out[18][4] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _5994_ (.RESET_B(net292),
    .D(_0044_),
    .Q(\s0.data_out[18][5] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _5995_ (.RESET_B(net291),
    .D(_0045_),
    .Q(\s0.data_out[18][6] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _5996_ (.RESET_B(net290),
    .D(_0046_),
    .Q(\s0.data_out[18][7] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _5997_ (.RESET_B(net289),
    .D(_0047_),
    .Q(\s0.shift_out[18] [0]),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _5998_ (.RESET_B(net288),
    .D(_0048_),
    .Q(\s0.genblk1[17].modules.bubble ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _5999_ (.RESET_B(net287),
    .D(net376),
    .Q(\s0.was_valid_out[17] [0]),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6000_ (.RESET_B(net285),
    .D(_0050_),
    .Q(\s0.valid_out[17] [0]),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _6001_ (.RESET_B(net284),
    .D(_0051_),
    .Q(\s0.data_out[17][0] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6002_ (.RESET_B(net283),
    .D(_0052_),
    .Q(\s0.data_out[17][1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6003_ (.RESET_B(net282),
    .D(_0053_),
    .Q(\s0.data_out[17][2] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6004_ (.RESET_B(net281),
    .D(_0054_),
    .Q(\s0.data_out[17][3] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6005_ (.RESET_B(net280),
    .D(_0055_),
    .Q(\s0.data_out[17][4] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _6006_ (.RESET_B(net279),
    .D(_0056_),
    .Q(\s0.data_out[17][5] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6007_ (.RESET_B(net278),
    .D(_0057_),
    .Q(\s0.data_out[17][6] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6008_ (.RESET_B(net277),
    .D(_0058_),
    .Q(\s0.data_out[17][7] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6009_ (.RESET_B(net276),
    .D(_0059_),
    .Q(\s0.shift_out[17] [0]),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6010_ (.RESET_B(net275),
    .D(_0060_),
    .Q(\s0.genblk1[16].modules.bubble ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6011_ (.RESET_B(net274),
    .D(net322),
    .Q(\s0.was_valid_out[16] [0]),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6012_ (.RESET_B(net272),
    .D(_0062_),
    .Q(\s0.valid_out[16] [0]),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6013_ (.RESET_B(net271),
    .D(_0063_),
    .Q(\s0.data_out[16][0] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6014_ (.RESET_B(net270),
    .D(_0064_),
    .Q(\s0.data_out[16][1] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6015_ (.RESET_B(net269),
    .D(_0065_),
    .Q(\s0.data_out[16][2] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6016_ (.RESET_B(net268),
    .D(_0066_),
    .Q(\s0.data_out[16][3] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6017_ (.RESET_B(net267),
    .D(_0067_),
    .Q(\s0.data_out[16][4] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6018_ (.RESET_B(net266),
    .D(_0068_),
    .Q(\s0.data_out[16][5] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6019_ (.RESET_B(net265),
    .D(_0069_),
    .Q(\s0.data_out[16][6] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6020_ (.RESET_B(net264),
    .D(_0070_),
    .Q(\s0.data_out[16][7] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6021_ (.RESET_B(net263),
    .D(_0071_),
    .Q(\s0.shift_out[16] [0]),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6022_ (.RESET_B(net262),
    .D(_0072_),
    .Q(\s0.genblk1[15].modules.bubble ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6023_ (.RESET_B(net261),
    .D(net382),
    .Q(\s0.was_valid_out[15] [0]),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6024_ (.RESET_B(net259),
    .D(_0074_),
    .Q(\s0.valid_out[15] [0]),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6025_ (.RESET_B(net258),
    .D(_0075_),
    .Q(\s0.data_out[15][0] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _6026_ (.RESET_B(net257),
    .D(_0076_),
    .Q(\s0.data_out[15][1] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _6027_ (.RESET_B(net256),
    .D(_0077_),
    .Q(\s0.data_out[15][2] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _6028_ (.RESET_B(net255),
    .D(_0078_),
    .Q(\s0.data_out[15][3] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _6029_ (.RESET_B(net254),
    .D(_0079_),
    .Q(\s0.data_out[15][4] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6030_ (.RESET_B(net253),
    .D(_0080_),
    .Q(\s0.data_out[15][5] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6031_ (.RESET_B(net252),
    .D(_0081_),
    .Q(\s0.data_out[15][6] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _6032_ (.RESET_B(net251),
    .D(_0082_),
    .Q(\s0.data_out[15][7] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6033_ (.RESET_B(net250),
    .D(_0083_),
    .Q(\s0.shift_out[15] [0]),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6034_ (.RESET_B(net249),
    .D(_0084_),
    .Q(\s0.genblk1[14].modules.bubble ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6035_ (.RESET_B(net248),
    .D(_0085_),
    .Q(\s0.was_valid_out[14] [0]),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6036_ (.RESET_B(net246),
    .D(_0086_),
    .Q(\s0.valid_out[14] [0]),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6037_ (.RESET_B(net245),
    .D(_0087_),
    .Q(\s0.data_out[14][0] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _6038_ (.RESET_B(net244),
    .D(_0088_),
    .Q(\s0.data_out[14][1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6039_ (.RESET_B(net243),
    .D(_0089_),
    .Q(\s0.data_out[14][2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6040_ (.RESET_B(net242),
    .D(_0090_),
    .Q(\s0.data_out[14][3] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6041_ (.RESET_B(net241),
    .D(_0091_),
    .Q(\s0.data_out[14][4] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6042_ (.RESET_B(net240),
    .D(_0092_),
    .Q(\s0.data_out[14][5] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6043_ (.RESET_B(net239),
    .D(_0093_),
    .Q(\s0.data_out[14][6] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _6044_ (.RESET_B(net238),
    .D(_0094_),
    .Q(\s0.data_out[14][7] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6045_ (.RESET_B(net237),
    .D(_0095_),
    .Q(\s0.shift_out[14] [0]),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6046_ (.RESET_B(net236),
    .D(_0096_),
    .Q(\s0.genblk1[13].modules.bubble ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6047_ (.RESET_B(net235),
    .D(net347),
    .Q(\s0.was_valid_out[13] [0]),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6048_ (.RESET_B(net233),
    .D(_0098_),
    .Q(\s0.valid_out[13] [0]),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6049_ (.RESET_B(net232),
    .D(_0099_),
    .Q(\s0.data_out[13][0] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6050_ (.RESET_B(net231),
    .D(_0100_),
    .Q(\s0.data_out[13][1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6051_ (.RESET_B(net230),
    .D(_0101_),
    .Q(\s0.data_out[13][2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6052_ (.RESET_B(net229),
    .D(_0102_),
    .Q(\s0.data_out[13][3] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6053_ (.RESET_B(net228),
    .D(_0103_),
    .Q(\s0.data_out[13][4] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6054_ (.RESET_B(net227),
    .D(_0104_),
    .Q(\s0.data_out[13][5] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6055_ (.RESET_B(net226),
    .D(_0105_),
    .Q(\s0.data_out[13][6] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6056_ (.RESET_B(net225),
    .D(_0106_),
    .Q(\s0.data_out[13][7] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6057_ (.RESET_B(net224),
    .D(_0107_),
    .Q(\s0.shift_out[13] [0]),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6058_ (.RESET_B(net223),
    .D(_0108_),
    .Q(\s0.genblk1[12].modules.bubble ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6059_ (.RESET_B(net222),
    .D(net409),
    .Q(\s0.was_valid_out[12] [0]),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6060_ (.RESET_B(net220),
    .D(_0110_),
    .Q(\s0.valid_out[12] [0]),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6061_ (.RESET_B(net219),
    .D(_0111_),
    .Q(\s0.data_out[12][0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6062_ (.RESET_B(net218),
    .D(_0112_),
    .Q(\s0.data_out[12][1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6063_ (.RESET_B(net217),
    .D(_0113_),
    .Q(\s0.data_out[12][2] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6064_ (.RESET_B(net216),
    .D(_0114_),
    .Q(\s0.data_out[12][3] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6065_ (.RESET_B(net215),
    .D(_0115_),
    .Q(\s0.data_out[12][4] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6066_ (.RESET_B(net214),
    .D(_0116_),
    .Q(\s0.data_out[12][5] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6067_ (.RESET_B(net213),
    .D(_0117_),
    .Q(\s0.data_out[12][6] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6068_ (.RESET_B(net212),
    .D(_0118_),
    .Q(\s0.data_out[12][7] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6069_ (.RESET_B(net211),
    .D(_0119_),
    .Q(\s0.shift_out[12] [0]),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6070_ (.RESET_B(net210),
    .D(_0120_),
    .Q(\s0.genblk1[11].modules.bubble ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6071_ (.RESET_B(net209),
    .D(_0121_),
    .Q(\s0.was_valid_out[11] [0]),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6072_ (.RESET_B(net207),
    .D(_0122_),
    .Q(\s0.valid_out[11] [0]),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6073_ (.RESET_B(net206),
    .D(_0123_),
    .Q(\s0.data_out[11][0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6074_ (.RESET_B(net205),
    .D(_0124_),
    .Q(\s0.data_out[11][1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6075_ (.RESET_B(net204),
    .D(_0125_),
    .Q(\s0.data_out[11][2] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _6076_ (.RESET_B(net203),
    .D(_0126_),
    .Q(\s0.data_out[11][3] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6077_ (.RESET_B(net202),
    .D(_0127_),
    .Q(\s0.data_out[11][4] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _6078_ (.RESET_B(net201),
    .D(_0128_),
    .Q(\s0.data_out[11][5] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6079_ (.RESET_B(net200),
    .D(_0129_),
    .Q(\s0.data_out[11][6] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _6080_ (.RESET_B(net199),
    .D(_0130_),
    .Q(\s0.data_out[11][7] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6081_ (.RESET_B(net198),
    .D(_0131_),
    .Q(\s0.shift_out[11] [0]),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6082_ (.RESET_B(net197),
    .D(_0132_),
    .Q(\s0.genblk1[10].modules.bubble ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6083_ (.RESET_B(net196),
    .D(net380),
    .Q(\s0.was_valid_out[10] [0]),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6084_ (.RESET_B(net194),
    .D(_0134_),
    .Q(\s0.valid_out[10] [0]),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _6085_ (.RESET_B(net193),
    .D(_0135_),
    .Q(\s0.data_out[10][0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6086_ (.RESET_B(net192),
    .D(_0136_),
    .Q(\s0.data_out[10][1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _6087_ (.RESET_B(net191),
    .D(_0137_),
    .Q(\s0.data_out[10][2] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _6088_ (.RESET_B(net190),
    .D(_0138_),
    .Q(\s0.data_out[10][3] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _6089_ (.RESET_B(net189),
    .D(_0139_),
    .Q(\s0.data_out[10][4] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _6090_ (.RESET_B(net188),
    .D(_0140_),
    .Q(\s0.data_out[10][5] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _6091_ (.RESET_B(net187),
    .D(_0141_),
    .Q(\s0.data_out[10][6] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _6092_ (.RESET_B(net186),
    .D(_0142_),
    .Q(\s0.data_out[10][7] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _6093_ (.RESET_B(net185),
    .D(_0143_),
    .Q(\s0.shift_out[10] [0]),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6094_ (.RESET_B(net184),
    .D(_0144_),
    .Q(\s0.data_new_delayed[0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6095_ (.RESET_B(net183),
    .D(_0145_),
    .Q(\s0.data_new_delayed[1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6096_ (.RESET_B(net182),
    .D(_0146_),
    .Q(\s0.data_new_delayed[2] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6097_ (.RESET_B(net181),
    .D(_0147_),
    .Q(\s0.data_new_delayed[3] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6098_ (.RESET_B(net180),
    .D(_0148_),
    .Q(\s0.data_new_delayed[4] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6099_ (.RESET_B(net179),
    .D(_0149_),
    .Q(\s0.data_new_delayed[5] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6100_ (.RESET_B(net178),
    .D(_0150_),
    .Q(\s0.data_new_delayed[6] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6101_ (.RESET_B(net177),
    .D(_0151_),
    .Q(\s0.data_new_delayed[7] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6102_ (.RESET_B(net176),
    .D(_0152_),
    .Q(\s0.was_valid_out[9] [0]),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6103_ (.RESET_B(net174),
    .D(_0153_),
    .Q(\s0.valid_out[9] [0]),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _6104_ (.RESET_B(net173),
    .D(_0154_),
    .Q(\s0.data_out[9][0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6105_ (.RESET_B(net172),
    .D(_0155_),
    .Q(\s0.data_out[9][1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6106_ (.RESET_B(net171),
    .D(_0156_),
    .Q(\s0.data_out[9][2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _6107_ (.RESET_B(net170),
    .D(_0157_),
    .Q(\s0.data_out[9][3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _6108_ (.RESET_B(net169),
    .D(_0158_),
    .Q(\s0.data_out[9][4] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _6109_ (.RESET_B(net168),
    .D(_0159_),
    .Q(\s0.data_out[9][5] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _6110_ (.RESET_B(net167),
    .D(_0160_),
    .Q(\s0.data_out[9][6] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _6111_ (.RESET_B(net166),
    .D(_0161_),
    .Q(\s0.data_out[9][7] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _6112_ (.RESET_B(net165),
    .D(_0162_),
    .Q(\s0.shift_out[9] [0]),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6113_ (.RESET_B(net164),
    .D(_0163_),
    .Q(\s0.genblk1[8].modules.bubble ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6114_ (.RESET_B(net163),
    .D(net399),
    .Q(\s0.was_valid_out[8] [0]),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6115_ (.RESET_B(net161),
    .D(_0165_),
    .Q(\s0.valid_out[8] [0]),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _6116_ (.RESET_B(net160),
    .D(_0166_),
    .Q(\s0.data_out[8][0] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6117_ (.RESET_B(net159),
    .D(_0167_),
    .Q(\s0.data_out[8][1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6118_ (.RESET_B(net158),
    .D(_0168_),
    .Q(\s0.data_out[8][2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _6119_ (.RESET_B(net157),
    .D(_0169_),
    .Q(\s0.data_out[8][3] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _6120_ (.RESET_B(net156),
    .D(_0170_),
    .Q(\s0.data_out[8][4] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _6121_ (.RESET_B(net155),
    .D(_0171_),
    .Q(\s0.data_out[8][5] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _6122_ (.RESET_B(net154),
    .D(_0172_),
    .Q(\s0.data_out[8][6] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _6123_ (.RESET_B(net153),
    .D(_0173_),
    .Q(\s0.data_out[8][7] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _6124_ (.RESET_B(net152),
    .D(_0174_),
    .Q(\s0.shift_out[8] [0]),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6125_ (.RESET_B(net151),
    .D(_0175_),
    .Q(\s0.genblk1[7].modules.bubble ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _6126_ (.RESET_B(net150),
    .D(net327),
    .Q(\s0.was_valid_out[7] [0]),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6127_ (.RESET_B(net148),
    .D(_0177_),
    .Q(\s0.valid_out[7] [0]),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _6128_ (.RESET_B(net147),
    .D(_0178_),
    .Q(\s0.data_out[7][0] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6129_ (.RESET_B(net146),
    .D(_0179_),
    .Q(\s0.data_out[7][1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6130_ (.RESET_B(net145),
    .D(_0180_),
    .Q(\s0.data_out[7][2] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _6131_ (.RESET_B(net144),
    .D(_0181_),
    .Q(\s0.data_out[7][3] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _6132_ (.RESET_B(net143),
    .D(_0182_),
    .Q(\s0.data_out[7][4] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _6133_ (.RESET_B(net142),
    .D(_0183_),
    .Q(\s0.data_out[7][5] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _6134_ (.RESET_B(net141),
    .D(_0184_),
    .Q(\s0.data_out[7][6] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _6135_ (.RESET_B(net140),
    .D(_0185_),
    .Q(\s0.data_out[7][7] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _6136_ (.RESET_B(net139),
    .D(_0186_),
    .Q(\s0.shift_out[7] [0]),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6137_ (.RESET_B(net138),
    .D(_0187_),
    .Q(\s0.genblk1[6].modules.bubble ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6138_ (.RESET_B(net137),
    .D(net466),
    .Q(\s0.was_valid_out[6] [0]),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6139_ (.RESET_B(net135),
    .D(_0189_),
    .Q(\s0.valid_out[6] [0]),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _6140_ (.RESET_B(net134),
    .D(_0190_),
    .Q(\s0.data_out[6][0] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6141_ (.RESET_B(net133),
    .D(_0191_),
    .Q(\s0.data_out[6][1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _6142_ (.RESET_B(net132),
    .D(_0192_),
    .Q(\s0.data_out[6][2] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _6143_ (.RESET_B(net131),
    .D(_0193_),
    .Q(\s0.data_out[6][3] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _6144_ (.RESET_B(net130),
    .D(_0194_),
    .Q(\s0.data_out[6][4] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _6145_ (.RESET_B(net129),
    .D(_0195_),
    .Q(\s0.data_out[6][5] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _6146_ (.RESET_B(net128),
    .D(_0196_),
    .Q(\s0.data_out[6][6] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _6147_ (.RESET_B(net127),
    .D(_0197_),
    .Q(\s0.data_out[6][7] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6148_ (.RESET_B(net126),
    .D(_0198_),
    .Q(\s0.shift_out[6] [0]),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6149_ (.RESET_B(net125),
    .D(_0199_),
    .Q(\s0.genblk1[5].modules.bubble ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6150_ (.RESET_B(net124),
    .D(net384),
    .Q(\s0.was_valid_out[5] [0]),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6151_ (.RESET_B(net122),
    .D(_0201_),
    .Q(\s0.valid_out[5] [0]),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _6152_ (.RESET_B(net121),
    .D(_0202_),
    .Q(\s0.data_out[5][0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _6153_ (.RESET_B(net120),
    .D(_0203_),
    .Q(\s0.data_out[5][1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _6154_ (.RESET_B(net119),
    .D(_0204_),
    .Q(\s0.data_out[5][2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _6155_ (.RESET_B(net118),
    .D(_0205_),
    .Q(\s0.data_out[5][3] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _6156_ (.RESET_B(net117),
    .D(_0206_),
    .Q(\s0.data_out[5][4] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _6157_ (.RESET_B(net116),
    .D(_0207_),
    .Q(\s0.data_out[5][5] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _6158_ (.RESET_B(net115),
    .D(_0208_),
    .Q(\s0.data_out[5][6] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _6159_ (.RESET_B(net114),
    .D(_0209_),
    .Q(\s0.data_out[5][7] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6160_ (.RESET_B(net113),
    .D(_0210_),
    .Q(\s0.shift_out[5] [0]),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6161_ (.RESET_B(net112),
    .D(_0211_),
    .Q(\s0.genblk1[4].modules.bubble ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6162_ (.RESET_B(net111),
    .D(_0212_),
    .Q(\s0.was_valid_out[4] [0]),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6163_ (.RESET_B(net109),
    .D(_0213_),
    .Q(\s0.valid_out[4] [0]),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _6164_ (.RESET_B(net108),
    .D(_0214_),
    .Q(\s0.data_out[4][0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _6165_ (.RESET_B(net107),
    .D(_0215_),
    .Q(\s0.data_out[4][1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _6166_ (.RESET_B(net106),
    .D(_0216_),
    .Q(\s0.data_out[4][2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _6167_ (.RESET_B(net105),
    .D(_0217_),
    .Q(\s0.data_out[4][3] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _6168_ (.RESET_B(net104),
    .D(_0218_),
    .Q(\s0.data_out[4][4] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _6169_ (.RESET_B(net103),
    .D(_0219_),
    .Q(\s0.data_out[4][5] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _6170_ (.RESET_B(net102),
    .D(_0220_),
    .Q(\s0.data_out[4][6] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _6171_ (.RESET_B(net101),
    .D(_0221_),
    .Q(\s0.data_out[4][7] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6172_ (.RESET_B(net100),
    .D(_0222_),
    .Q(\s0.shift_out[4] [0]),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6173_ (.RESET_B(net99),
    .D(_0223_),
    .Q(\s0.genblk1[3].modules.bubble ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6174_ (.RESET_B(net98),
    .D(net320),
    .Q(\s0.was_valid_out[3] [0]),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6175_ (.RESET_B(net96),
    .D(_0225_),
    .Q(\s0.valid_out[3] [0]),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _6176_ (.RESET_B(net95),
    .D(_0226_),
    .Q(\s0.data_out[3][0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _6177_ (.RESET_B(net94),
    .D(_0227_),
    .Q(\s0.data_out[3][1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _6178_ (.RESET_B(net93),
    .D(_0228_),
    .Q(\s0.data_out[3][2] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _6179_ (.RESET_B(net92),
    .D(_0229_),
    .Q(\s0.data_out[3][3] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _6180_ (.RESET_B(net91),
    .D(_0230_),
    .Q(\s0.data_out[3][4] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _6181_ (.RESET_B(net90),
    .D(_0231_),
    .Q(\s0.data_out[3][5] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _6182_ (.RESET_B(net89),
    .D(_0232_),
    .Q(\s0.data_out[3][6] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _6183_ (.RESET_B(net88),
    .D(_0233_),
    .Q(\s0.data_out[3][7] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6184_ (.RESET_B(net87),
    .D(_0234_),
    .Q(\s0.shift_out[3] [0]),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6185_ (.RESET_B(net86),
    .D(_0235_),
    .Q(\s0.genblk1[2].modules.bubble ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6186_ (.RESET_B(net85),
    .D(_0236_),
    .Q(\s0.was_valid_out[2] [0]),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6187_ (.RESET_B(net83),
    .D(_0237_),
    .Q(\s0.valid_out[2] [0]),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6188_ (.RESET_B(net82),
    .D(_0238_),
    .Q(\s0.data_out[2][0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _6189_ (.RESET_B(net81),
    .D(_0239_),
    .Q(\s0.data_out[2][1] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _6190_ (.RESET_B(net80),
    .D(_0240_),
    .Q(\s0.data_out[2][2] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _6191_ (.RESET_B(net79),
    .D(_0241_),
    .Q(\s0.data_out[2][3] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6192_ (.RESET_B(net78),
    .D(_0242_),
    .Q(\s0.data_out[2][4] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6193_ (.RESET_B(net77),
    .D(_0243_),
    .Q(\s0.data_out[2][5] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _6194_ (.RESET_B(net76),
    .D(_0244_),
    .Q(\s0.data_out[2][6] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _6195_ (.RESET_B(net75),
    .D(_0245_),
    .Q(\s0.data_out[2][7] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _6196_ (.RESET_B(net74),
    .D(_0246_),
    .Q(\s0.shift_out[2] [0]),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6197_ (.RESET_B(net73),
    .D(_0247_),
    .Q(\s0.genblk1[21].modules.bubble ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6198_ (.RESET_B(net72),
    .D(net329),
    .Q(\s0.was_valid_out[1] [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6199_ (.RESET_B(net70),
    .D(_0249_),
    .Q(\s0.valid_out[1] [0]),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _6200_ (.RESET_B(net69),
    .D(_0250_),
    .Q(\s0.data_out[1][0] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _6201_ (.RESET_B(net68),
    .D(_0251_),
    .Q(\s0.data_out[1][1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _6202_ (.RESET_B(net66),
    .D(_0252_),
    .Q(\s0.data_out[1][2] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6203_ (.RESET_B(net53),
    .D(_0253_),
    .Q(\s0.data_out[1][3] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6204_ (.RESET_B(net40),
    .D(_0254_),
    .Q(\s0.data_out[1][4] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6205_ (.RESET_B(net27),
    .D(_0255_),
    .Q(\s0.data_out[1][5] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _6206_ (.RESET_B(net286),
    .D(_0256_),
    .Q(\s0.data_out[1][6] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _6207_ (.RESET_B(net273),
    .D(_0257_),
    .Q(\s0.data_out[1][7] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _6208_ (.RESET_B(net260),
    .D(_0258_),
    .Q(\s0.shift_out[1] [0]),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6209_ (.RESET_B(net247),
    .D(_0259_),
    .Q(\s0.genblk1[19].modules.bubble ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6210_ (.RESET_B(net234),
    .D(_0260_),
    .Q(\s0.was_valid_out[0] [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6211_ (.RESET_B(net208),
    .D(_0261_),
    .Q(\s0.valid_out[0] [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _6212_ (.RESET_B(net195),
    .D(_0262_),
    .Q(\s0.data_out[0][0] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _6213_ (.RESET_B(net175),
    .D(_0263_),
    .Q(\s0.data_out[0][1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6214_ (.RESET_B(net162),
    .D(_0264_),
    .Q(\s0.data_out[0][2] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6215_ (.RESET_B(net149),
    .D(_0265_),
    .Q(\s0.data_out[0][3] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _6216_ (.RESET_B(net136),
    .D(_0266_),
    .Q(\s0.data_out[0][4] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6217_ (.RESET_B(net123),
    .D(_0267_),
    .Q(\s0.data_out[0][5] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _6218_ (.RESET_B(net110),
    .D(_0268_),
    .Q(\s0.data_out[0][6] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6219_ (.RESET_B(net97),
    .D(_0269_),
    .Q(\s0.data_out[0][7] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6220_ (.RESET_B(net84),
    .D(_0270_),
    .Q(\s0.shift_out[0] [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6221_ (.RESET_B(net71),
    .D(_0271_),
    .Q(\s0.genblk1[9].modules.bubble ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_tiehi _5990__24 (.L_HI(net24));
 sg13g2_tiehi _5989__25 (.L_HI(net25));
 sg13g2_tiehi _5988__26 (.L_HI(net26));
 sg13g2_tiehi _6205__27 (.L_HI(net27));
 sg13g2_tiehi _5987__28 (.L_HI(net28));
 sg13g2_tiehi _5986__29 (.L_HI(net29));
 sg13g2_tiehi _5985__30 (.L_HI(net30));
 sg13g2_tiehi _5984__31 (.L_HI(net31));
 sg13g2_tiehi _5983__32 (.L_HI(net32));
 sg13g2_tiehi _5982__33 (.L_HI(net33));
 sg13g2_tiehi _5981__34 (.L_HI(net34));
 sg13g2_tiehi _5980__35 (.L_HI(net35));
 sg13g2_tiehi _5979__36 (.L_HI(net36));
 sg13g2_tiehi _5978__37 (.L_HI(net37));
 sg13g2_tiehi _5977__38 (.L_HI(net38));
 sg13g2_tiehi _5976__39 (.L_HI(net39));
 sg13g2_tiehi _6204__40 (.L_HI(net40));
 sg13g2_tiehi _5975__41 (.L_HI(net41));
 sg13g2_tiehi _5974__42 (.L_HI(net42));
 sg13g2_tiehi _5973__43 (.L_HI(net43));
 sg13g2_tiehi _5972__44 (.L_HI(net44));
 sg13g2_tiehi _5971__45 (.L_HI(net45));
 sg13g2_tiehi _5970__46 (.L_HI(net46));
 sg13g2_tiehi _5969__47 (.L_HI(net47));
 sg13g2_tiehi _5968__48 (.L_HI(net48));
 sg13g2_tiehi _5967__49 (.L_HI(net49));
 sg13g2_tiehi _5966__50 (.L_HI(net50));
 sg13g2_tiehi _5965__51 (.L_HI(net51));
 sg13g2_tiehi _5964__52 (.L_HI(net52));
 sg13g2_tiehi _6203__53 (.L_HI(net53));
 sg13g2_tiehi _5963__54 (.L_HI(net54));
 sg13g2_tiehi _5962__55 (.L_HI(net55));
 sg13g2_tiehi _5961__56 (.L_HI(net56));
 sg13g2_tiehi _5960__57 (.L_HI(net57));
 sg13g2_tiehi _5959__58 (.L_HI(net58));
 sg13g2_tiehi _5958__59 (.L_HI(net59));
 sg13g2_tiehi _5957__60 (.L_HI(net60));
 sg13g2_tiehi _5956__61 (.L_HI(net61));
 sg13g2_tiehi _5955__62 (.L_HI(net62));
 sg13g2_tiehi _5954__63 (.L_HI(net63));
 sg13g2_tiehi _5953__64 (.L_HI(net64));
 sg13g2_tiehi _5952__65 (.L_HI(net65));
 sg13g2_tiehi _6202__66 (.L_HI(net66));
 sg13g2_tiehi _5951__67 (.L_HI(net67));
 sg13g2_tiehi _6201__68 (.L_HI(net68));
 sg13g2_tiehi _6200__69 (.L_HI(net69));
 sg13g2_tiehi _6199__70 (.L_HI(net70));
 sg13g2_tiehi _6221__71 (.L_HI(net71));
 sg13g2_tiehi _6198__72 (.L_HI(net72));
 sg13g2_tiehi _6197__73 (.L_HI(net73));
 sg13g2_tiehi _6196__74 (.L_HI(net74));
 sg13g2_tiehi _6195__75 (.L_HI(net75));
 sg13g2_tiehi _6194__76 (.L_HI(net76));
 sg13g2_tiehi _6193__77 (.L_HI(net77));
 sg13g2_tiehi _6192__78 (.L_HI(net78));
 sg13g2_tiehi _6191__79 (.L_HI(net79));
 sg13g2_tiehi _6190__80 (.L_HI(net80));
 sg13g2_tiehi _6189__81 (.L_HI(net81));
 sg13g2_tiehi _6188__82 (.L_HI(net82));
 sg13g2_tiehi _6187__83 (.L_HI(net83));
 sg13g2_tiehi _6220__84 (.L_HI(net84));
 sg13g2_tiehi _6186__85 (.L_HI(net85));
 sg13g2_tiehi _6185__86 (.L_HI(net86));
 sg13g2_tiehi _6184__87 (.L_HI(net87));
 sg13g2_tiehi _6183__88 (.L_HI(net88));
 sg13g2_tiehi _6182__89 (.L_HI(net89));
 sg13g2_tiehi _6181__90 (.L_HI(net90));
 sg13g2_tiehi _6180__91 (.L_HI(net91));
 sg13g2_tiehi _6179__92 (.L_HI(net92));
 sg13g2_tiehi _6178__93 (.L_HI(net93));
 sg13g2_tiehi _6177__94 (.L_HI(net94));
 sg13g2_tiehi _6176__95 (.L_HI(net95));
 sg13g2_tiehi _6175__96 (.L_HI(net96));
 sg13g2_tiehi _6219__97 (.L_HI(net97));
 sg13g2_tiehi _6174__98 (.L_HI(net98));
 sg13g2_tiehi _6173__99 (.L_HI(net99));
 sg13g2_tiehi _6172__100 (.L_HI(net100));
 sg13g2_tiehi _6171__101 (.L_HI(net101));
 sg13g2_tiehi _6170__102 (.L_HI(net102));
 sg13g2_tiehi _6169__103 (.L_HI(net103));
 sg13g2_tiehi _6168__104 (.L_HI(net104));
 sg13g2_tiehi _6167__105 (.L_HI(net105));
 sg13g2_tiehi _6166__106 (.L_HI(net106));
 sg13g2_tiehi _6165__107 (.L_HI(net107));
 sg13g2_tiehi _6164__108 (.L_HI(net108));
 sg13g2_tiehi _6163__109 (.L_HI(net109));
 sg13g2_tiehi _6218__110 (.L_HI(net110));
 sg13g2_tiehi _6162__111 (.L_HI(net111));
 sg13g2_tiehi _6161__112 (.L_HI(net112));
 sg13g2_tiehi _6160__113 (.L_HI(net113));
 sg13g2_tiehi _6159__114 (.L_HI(net114));
 sg13g2_tiehi _6158__115 (.L_HI(net115));
 sg13g2_tiehi _6157__116 (.L_HI(net116));
 sg13g2_tiehi _6156__117 (.L_HI(net117));
 sg13g2_tiehi _6155__118 (.L_HI(net118));
 sg13g2_tiehi _6154__119 (.L_HI(net119));
 sg13g2_tiehi _6153__120 (.L_HI(net120));
 sg13g2_tiehi _6152__121 (.L_HI(net121));
 sg13g2_tiehi _6151__122 (.L_HI(net122));
 sg13g2_tiehi _6217__123 (.L_HI(net123));
 sg13g2_tiehi _6150__124 (.L_HI(net124));
 sg13g2_tiehi _6149__125 (.L_HI(net125));
 sg13g2_tiehi _6148__126 (.L_HI(net126));
 sg13g2_tiehi _6147__127 (.L_HI(net127));
 sg13g2_tiehi _6146__128 (.L_HI(net128));
 sg13g2_tiehi _6145__129 (.L_HI(net129));
 sg13g2_tiehi _6144__130 (.L_HI(net130));
 sg13g2_tiehi _6143__131 (.L_HI(net131));
 sg13g2_tiehi _6142__132 (.L_HI(net132));
 sg13g2_tiehi _6141__133 (.L_HI(net133));
 sg13g2_tiehi _6140__134 (.L_HI(net134));
 sg13g2_tiehi _6139__135 (.L_HI(net135));
 sg13g2_tiehi _6216__136 (.L_HI(net136));
 sg13g2_tiehi _6138__137 (.L_HI(net137));
 sg13g2_tiehi _6137__138 (.L_HI(net138));
 sg13g2_tiehi _6136__139 (.L_HI(net139));
 sg13g2_tiehi _6135__140 (.L_HI(net140));
 sg13g2_tiehi _6134__141 (.L_HI(net141));
 sg13g2_tiehi _6133__142 (.L_HI(net142));
 sg13g2_tiehi _6132__143 (.L_HI(net143));
 sg13g2_tiehi _6131__144 (.L_HI(net144));
 sg13g2_tiehi _6130__145 (.L_HI(net145));
 sg13g2_tiehi _6129__146 (.L_HI(net146));
 sg13g2_tiehi _6128__147 (.L_HI(net147));
 sg13g2_tiehi _6127__148 (.L_HI(net148));
 sg13g2_tiehi _6215__149 (.L_HI(net149));
 sg13g2_tiehi _6126__150 (.L_HI(net150));
 sg13g2_tiehi _6125__151 (.L_HI(net151));
 sg13g2_tiehi _6124__152 (.L_HI(net152));
 sg13g2_tiehi _6123__153 (.L_HI(net153));
 sg13g2_tiehi _6122__154 (.L_HI(net154));
 sg13g2_tiehi _6121__155 (.L_HI(net155));
 sg13g2_tiehi _6120__156 (.L_HI(net156));
 sg13g2_tiehi _6119__157 (.L_HI(net157));
 sg13g2_tiehi _6118__158 (.L_HI(net158));
 sg13g2_tiehi _6117__159 (.L_HI(net159));
 sg13g2_tiehi _6116__160 (.L_HI(net160));
 sg13g2_tiehi _6115__161 (.L_HI(net161));
 sg13g2_tiehi _6214__162 (.L_HI(net162));
 sg13g2_tiehi _6114__163 (.L_HI(net163));
 sg13g2_tiehi _6113__164 (.L_HI(net164));
 sg13g2_tiehi _6112__165 (.L_HI(net165));
 sg13g2_tiehi _6111__166 (.L_HI(net166));
 sg13g2_tiehi _6110__167 (.L_HI(net167));
 sg13g2_tiehi _6109__168 (.L_HI(net168));
 sg13g2_tiehi _6108__169 (.L_HI(net169));
 sg13g2_tiehi _6107__170 (.L_HI(net170));
 sg13g2_tiehi _6106__171 (.L_HI(net171));
 sg13g2_tiehi _6105__172 (.L_HI(net172));
 sg13g2_tiehi _6104__173 (.L_HI(net173));
 sg13g2_tiehi _6103__174 (.L_HI(net174));
 sg13g2_tiehi _6213__175 (.L_HI(net175));
 sg13g2_tiehi _6102__176 (.L_HI(net176));
 sg13g2_tiehi _6101__177 (.L_HI(net177));
 sg13g2_tiehi _6100__178 (.L_HI(net178));
 sg13g2_tiehi _6099__179 (.L_HI(net179));
 sg13g2_tiehi _6098__180 (.L_HI(net180));
 sg13g2_tiehi _6097__181 (.L_HI(net181));
 sg13g2_tiehi _6096__182 (.L_HI(net182));
 sg13g2_tiehi _6095__183 (.L_HI(net183));
 sg13g2_tiehi _6094__184 (.L_HI(net184));
 sg13g2_tiehi _6093__185 (.L_HI(net185));
 sg13g2_tiehi _6092__186 (.L_HI(net186));
 sg13g2_tiehi _6091__187 (.L_HI(net187));
 sg13g2_tiehi _6090__188 (.L_HI(net188));
 sg13g2_tiehi _6089__189 (.L_HI(net189));
 sg13g2_tiehi _6088__190 (.L_HI(net190));
 sg13g2_tiehi _6087__191 (.L_HI(net191));
 sg13g2_tiehi _6086__192 (.L_HI(net192));
 sg13g2_tiehi _6085__193 (.L_HI(net193));
 sg13g2_tiehi _6084__194 (.L_HI(net194));
 sg13g2_tiehi _6212__195 (.L_HI(net195));
 sg13g2_tiehi _6083__196 (.L_HI(net196));
 sg13g2_tiehi _6082__197 (.L_HI(net197));
 sg13g2_tiehi _6081__198 (.L_HI(net198));
 sg13g2_tiehi _6080__199 (.L_HI(net199));
 sg13g2_tiehi _6079__200 (.L_HI(net200));
 sg13g2_tiehi _6078__201 (.L_HI(net201));
 sg13g2_tiehi _6077__202 (.L_HI(net202));
 sg13g2_tiehi _6076__203 (.L_HI(net203));
 sg13g2_tiehi _6075__204 (.L_HI(net204));
 sg13g2_tiehi _6074__205 (.L_HI(net205));
 sg13g2_tiehi _6073__206 (.L_HI(net206));
 sg13g2_tiehi _6072__207 (.L_HI(net207));
 sg13g2_tiehi _6211__208 (.L_HI(net208));
 sg13g2_tiehi _6071__209 (.L_HI(net209));
 sg13g2_tiehi _6070__210 (.L_HI(net210));
 sg13g2_tiehi _6069__211 (.L_HI(net211));
 sg13g2_tiehi _6068__212 (.L_HI(net212));
 sg13g2_tiehi _6067__213 (.L_HI(net213));
 sg13g2_tiehi _6066__214 (.L_HI(net214));
 sg13g2_tiehi _6065__215 (.L_HI(net215));
 sg13g2_tiehi _6064__216 (.L_HI(net216));
 sg13g2_tiehi _6063__217 (.L_HI(net217));
 sg13g2_tiehi _6062__218 (.L_HI(net218));
 sg13g2_tiehi _6061__219 (.L_HI(net219));
 sg13g2_tiehi _6060__220 (.L_HI(net220));
 sg13g2_tiehi _5950__221 (.L_HI(net221));
 sg13g2_tiehi _6059__222 (.L_HI(net222));
 sg13g2_tiehi _6058__223 (.L_HI(net223));
 sg13g2_tiehi _6057__224 (.L_HI(net224));
 sg13g2_tiehi _6056__225 (.L_HI(net225));
 sg13g2_tiehi _6055__226 (.L_HI(net226));
 sg13g2_tiehi _6054__227 (.L_HI(net227));
 sg13g2_tiehi _6053__228 (.L_HI(net228));
 sg13g2_tiehi _6052__229 (.L_HI(net229));
 sg13g2_tiehi _6051__230 (.L_HI(net230));
 sg13g2_tiehi _6050__231 (.L_HI(net231));
 sg13g2_tiehi _6049__232 (.L_HI(net232));
 sg13g2_tiehi _6048__233 (.L_HI(net233));
 sg13g2_tiehi _6210__234 (.L_HI(net234));
 sg13g2_tiehi _6047__235 (.L_HI(net235));
 sg13g2_tiehi _6046__236 (.L_HI(net236));
 sg13g2_tiehi _6045__237 (.L_HI(net237));
 sg13g2_tiehi _6044__238 (.L_HI(net238));
 sg13g2_tiehi _6043__239 (.L_HI(net239));
 sg13g2_tiehi _6042__240 (.L_HI(net240));
 sg13g2_tiehi _6041__241 (.L_HI(net241));
 sg13g2_tiehi _6040__242 (.L_HI(net242));
 sg13g2_tiehi _6039__243 (.L_HI(net243));
 sg13g2_tiehi _6038__244 (.L_HI(net244));
 sg13g2_tiehi _6037__245 (.L_HI(net245));
 sg13g2_tiehi _6036__246 (.L_HI(net246));
 sg13g2_tiehi _6209__247 (.L_HI(net247));
 sg13g2_tiehi _6035__248 (.L_HI(net248));
 sg13g2_tiehi _6034__249 (.L_HI(net249));
 sg13g2_tiehi _6033__250 (.L_HI(net250));
 sg13g2_tiehi _6032__251 (.L_HI(net251));
 sg13g2_tiehi _6031__252 (.L_HI(net252));
 sg13g2_tiehi _6030__253 (.L_HI(net253));
 sg13g2_tiehi _6029__254 (.L_HI(net254));
 sg13g2_tiehi _6028__255 (.L_HI(net255));
 sg13g2_tiehi _6027__256 (.L_HI(net256));
 sg13g2_tiehi _6026__257 (.L_HI(net257));
 sg13g2_tiehi _6025__258 (.L_HI(net258));
 sg13g2_tiehi _6024__259 (.L_HI(net259));
 sg13g2_tiehi _6208__260 (.L_HI(net260));
 sg13g2_tiehi _6023__261 (.L_HI(net261));
 sg13g2_tiehi _6022__262 (.L_HI(net262));
 sg13g2_tiehi _6021__263 (.L_HI(net263));
 sg13g2_tiehi _6020__264 (.L_HI(net264));
 sg13g2_tiehi _6019__265 (.L_HI(net265));
 sg13g2_tiehi _6018__266 (.L_HI(net266));
 sg13g2_tiehi _6017__267 (.L_HI(net267));
 sg13g2_tiehi _6016__268 (.L_HI(net268));
 sg13g2_tiehi _6015__269 (.L_HI(net269));
 sg13g2_tiehi _6014__270 (.L_HI(net270));
 sg13g2_tiehi _6013__271 (.L_HI(net271));
 sg13g2_tiehi _6012__272 (.L_HI(net272));
 sg13g2_tiehi _6207__273 (.L_HI(net273));
 sg13g2_tiehi _6011__274 (.L_HI(net274));
 sg13g2_tiehi _6010__275 (.L_HI(net275));
 sg13g2_tiehi _6009__276 (.L_HI(net276));
 sg13g2_tiehi _6008__277 (.L_HI(net277));
 sg13g2_tiehi _6007__278 (.L_HI(net278));
 sg13g2_tiehi _6006__279 (.L_HI(net279));
 sg13g2_tiehi _6005__280 (.L_HI(net280));
 sg13g2_tiehi _6004__281 (.L_HI(net281));
 sg13g2_tiehi _6003__282 (.L_HI(net282));
 sg13g2_tiehi _6002__283 (.L_HI(net283));
 sg13g2_tiehi _6001__284 (.L_HI(net284));
 sg13g2_tiehi _6000__285 (.L_HI(net285));
 sg13g2_tiehi _6206__286 (.L_HI(net286));
 sg13g2_tiehi _5999__287 (.L_HI(net287));
 sg13g2_tiehi _5998__288 (.L_HI(net288));
 sg13g2_tiehi _5997__289 (.L_HI(net289));
 sg13g2_tiehi _5996__290 (.L_HI(net290));
 sg13g2_tiehi _5995__291 (.L_HI(net291));
 sg13g2_tiehi _5994__292 (.L_HI(net292));
 sg13g2_tiehi _5993__293 (.L_HI(net293));
 sg13g2_tiehi _5992__294 (.L_HI(net294));
 sg13g2_tiehi heichips25_top_sorter_295 (.L_HI(net295));
 sg13g2_tiehi heichips25_top_sorter_296 (.L_HI(net296));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo heichips25_top_sorter_11 (.L_LO(net11));
 sg13g2_tielo heichips25_top_sorter_12 (.L_LO(net12));
 sg13g2_tielo heichips25_top_sorter_13 (.L_LO(net13));
 sg13g2_tielo heichips25_top_sorter_14 (.L_LO(net14));
 sg13g2_tielo heichips25_top_sorter_15 (.L_LO(net15));
 sg13g2_tielo heichips25_top_sorter_16 (.L_LO(net16));
 sg13g2_tielo heichips25_top_sorter_17 (.L_LO(net17));
 sg13g2_tielo heichips25_top_sorter_18 (.L_LO(net18));
 sg13g2_tielo heichips25_top_sorter_19 (.L_LO(net19));
 sg13g2_tielo heichips25_top_sorter_20 (.L_LO(net20));
 sg13g2_tielo heichips25_top_sorter_21 (.L_LO(net21));
 sg13g2_tielo heichips25_top_sorter_22 (.L_LO(net22));
 sg13g2_tiehi _5991__23 (.L_HI(net23));
 sg13g2_buf_1 _6509_ (.A(\s0.was_valid_out[21] [0]),
    .X(net1));
 sg13g2_buf_8 fanout912 (.A(net913),
    .X(net912));
 sg13g2_buf_8 fanout913 (.A(_2494_),
    .X(net913));
 sg13g2_buf_8 fanout914 (.A(_2471_),
    .X(net914));
 sg13g2_buf_8 fanout915 (.A(_2470_),
    .X(net915));
 sg13g2_buf_8 fanout916 (.A(_2469_),
    .X(net916));
 sg13g2_buf_8 fanout917 (.A(_2468_),
    .X(net917));
 sg13g2_buf_8 fanout918 (.A(_2467_),
    .X(net918));
 sg13g2_buf_8 fanout919 (.A(_2466_),
    .X(net919));
 sg13g2_buf_1 fanout920 (.A(_2466_),
    .X(net920));
 sg13g2_buf_8 fanout921 (.A(_2464_),
    .X(net921));
 sg13g2_buf_8 fanout922 (.A(_2463_),
    .X(net922));
 sg13g2_buf_1 fanout923 (.A(_2463_),
    .X(net923));
 sg13g2_buf_8 fanout924 (.A(_2462_),
    .X(net924));
 sg13g2_buf_8 fanout925 (.A(_2461_),
    .X(net925));
 sg13g2_buf_8 fanout926 (.A(_2460_),
    .X(net926));
 sg13g2_buf_1 fanout927 (.A(_2460_),
    .X(net927));
 sg13g2_buf_8 fanout928 (.A(_2459_),
    .X(net928));
 sg13g2_buf_1 fanout929 (.A(_2459_),
    .X(net929));
 sg13g2_buf_8 fanout930 (.A(_2458_),
    .X(net930));
 sg13g2_buf_8 fanout931 (.A(_2456_),
    .X(net931));
 sg13g2_buf_8 fanout932 (.A(_2455_),
    .X(net932));
 sg13g2_buf_1 fanout933 (.A(_2455_),
    .X(net933));
 sg13g2_buf_8 fanout934 (.A(_2454_),
    .X(net934));
 sg13g2_buf_8 fanout935 (.A(_2453_),
    .X(net935));
 sg13g2_buf_1 fanout936 (.A(_2453_),
    .X(net936));
 sg13g2_buf_8 fanout937 (.A(_2452_),
    .X(net937));
 sg13g2_buf_8 fanout938 (.A(_2451_),
    .X(net938));
 sg13g2_buf_8 fanout939 (.A(_2448_),
    .X(net939));
 sg13g2_buf_2 fanout940 (.A(net941),
    .X(net940));
 sg13g2_buf_2 fanout941 (.A(net942),
    .X(net941));
 sg13g2_buf_8 fanout942 (.A(net945),
    .X(net942));
 sg13g2_buf_8 fanout943 (.A(net944),
    .X(net943));
 sg13g2_buf_8 fanout944 (.A(net945),
    .X(net944));
 sg13g2_buf_8 fanout945 (.A(net354),
    .X(net945));
 sg13g2_buf_8 fanout946 (.A(net948),
    .X(net946));
 sg13g2_buf_8 fanout947 (.A(net948),
    .X(net947));
 sg13g2_buf_8 fanout948 (.A(\s0.valid_out[0] [0]),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(net950),
    .X(net949));
 sg13g2_buf_8 fanout950 (.A(net951),
    .X(net950));
 sg13g2_buf_8 fanout951 (.A(\s0.shift_out[1] [0]),
    .X(net951));
 sg13g2_buf_8 fanout952 (.A(net954),
    .X(net952));
 sg13g2_buf_8 fanout953 (.A(net954),
    .X(net953));
 sg13g2_buf_8 fanout954 (.A(\s0.shift_out[1] [0]),
    .X(net954));
 sg13g2_buf_8 fanout955 (.A(net958),
    .X(net955));
 sg13g2_buf_8 fanout956 (.A(net958),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(net958),
    .X(net957));
 sg13g2_buf_8 fanout958 (.A(\s0.valid_out[1] [0]),
    .X(net958));
 sg13g2_buf_8 fanout959 (.A(net960),
    .X(net959));
 sg13g2_buf_8 fanout960 (.A(\s0.shift_out[2] [0]),
    .X(net960));
 sg13g2_buf_8 fanout961 (.A(\s0.shift_out[2] [0]),
    .X(net961));
 sg13g2_buf_8 fanout962 (.A(net964),
    .X(net962));
 sg13g2_buf_8 fanout963 (.A(net964),
    .X(net963));
 sg13g2_buf_8 fanout964 (.A(\s0.shift_out[2] [0]),
    .X(net964));
 sg13g2_buf_8 fanout965 (.A(net968),
    .X(net965));
 sg13g2_buf_8 fanout966 (.A(net968),
    .X(net966));
 sg13g2_buf_1 fanout967 (.A(net968),
    .X(net967));
 sg13g2_buf_8 fanout968 (.A(\s0.valid_out[2] [0]),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(net970),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(net975),
    .X(net970));
 sg13g2_buf_8 fanout971 (.A(net975),
    .X(net971));
 sg13g2_buf_8 fanout972 (.A(net974),
    .X(net972));
 sg13g2_buf_8 fanout973 (.A(net975),
    .X(net973));
 sg13g2_buf_1 fanout974 (.A(net975),
    .X(net974));
 sg13g2_buf_8 fanout975 (.A(\s0.shift_out[3] [0]),
    .X(net975));
 sg13g2_buf_8 fanout976 (.A(net979),
    .X(net976));
 sg13g2_buf_8 fanout977 (.A(net979),
    .X(net977));
 sg13g2_buf_1 fanout978 (.A(net979),
    .X(net978));
 sg13g2_buf_8 fanout979 (.A(\s0.valid_out[3] [0]),
    .X(net979));
 sg13g2_buf_8 fanout980 (.A(net986),
    .X(net980));
 sg13g2_buf_8 fanout981 (.A(net982),
    .X(net981));
 sg13g2_buf_8 fanout982 (.A(net986),
    .X(net982));
 sg13g2_buf_8 fanout983 (.A(net985),
    .X(net983));
 sg13g2_buf_8 fanout984 (.A(net985),
    .X(net984));
 sg13g2_buf_8 fanout985 (.A(net986),
    .X(net985));
 sg13g2_buf_8 fanout986 (.A(\s0.shift_out[4] [0]),
    .X(net986));
 sg13g2_buf_8 fanout987 (.A(net989),
    .X(net987));
 sg13g2_buf_8 fanout988 (.A(net989),
    .X(net988));
 sg13g2_buf_8 fanout989 (.A(\s0.valid_out[4] [0]),
    .X(net989));
 sg13g2_buf_8 fanout990 (.A(net993),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(net992),
    .X(net991));
 sg13g2_buf_8 fanout992 (.A(net993),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(\s0.shift_out[5] [0]),
    .X(net993));
 sg13g2_buf_8 fanout994 (.A(net996),
    .X(net994));
 sg13g2_buf_8 fanout995 (.A(net996),
    .X(net995));
 sg13g2_buf_8 fanout996 (.A(\s0.shift_out[5] [0]),
    .X(net996));
 sg13g2_buf_8 fanout997 (.A(net999),
    .X(net997));
 sg13g2_buf_8 fanout998 (.A(net999),
    .X(net998));
 sg13g2_buf_8 fanout999 (.A(\s0.valid_out[5] [0]),
    .X(net999));
 sg13g2_buf_8 fanout1000 (.A(net1003),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(net1002),
    .X(net1001));
 sg13g2_buf_1 fanout1002 (.A(net1003),
    .X(net1002));
 sg13g2_buf_1 fanout1003 (.A(\s0.shift_out[6] [0]),
    .X(net1003));
 sg13g2_buf_8 fanout1004 (.A(net1007),
    .X(net1004));
 sg13g2_buf_8 fanout1005 (.A(net1007),
    .X(net1005));
 sg13g2_buf_1 fanout1006 (.A(net1007),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(\s0.shift_out[6] [0]),
    .X(net1007));
 sg13g2_buf_8 fanout1008 (.A(net1011),
    .X(net1008));
 sg13g2_buf_8 fanout1009 (.A(net1011),
    .X(net1009));
 sg13g2_buf_2 fanout1010 (.A(net1011),
    .X(net1010));
 sg13g2_buf_8 fanout1011 (.A(\s0.valid_out[6] [0]),
    .X(net1011));
 sg13g2_buf_8 fanout1012 (.A(net340),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(net1014),
    .X(net1013));
 sg13g2_buf_8 fanout1014 (.A(\s0.shift_out[7] [0]),
    .X(net1014));
 sg13g2_buf_8 fanout1015 (.A(net1018),
    .X(net1015));
 sg13g2_buf_8 fanout1016 (.A(net1018),
    .X(net1016));
 sg13g2_buf_1 fanout1017 (.A(net1018),
    .X(net1017));
 sg13g2_buf_8 fanout1018 (.A(net339),
    .X(net1018));
 sg13g2_buf_8 fanout1019 (.A(net1022),
    .X(net1019));
 sg13g2_buf_8 fanout1020 (.A(net1021),
    .X(net1020));
 sg13g2_buf_8 fanout1021 (.A(net1022),
    .X(net1021));
 sg13g2_buf_8 fanout1022 (.A(\s0.valid_out[7] [0]),
    .X(net1022));
 sg13g2_buf_8 fanout1023 (.A(net1026),
    .X(net1023));
 sg13g2_buf_1 fanout1024 (.A(net1026),
    .X(net1024));
 sg13g2_buf_8 fanout1025 (.A(net1026),
    .X(net1025));
 sg13g2_buf_8 fanout1026 (.A(\s0.shift_out[8] [0]),
    .X(net1026));
 sg13g2_buf_8 fanout1027 (.A(net1029),
    .X(net1027));
 sg13g2_buf_1 fanout1028 (.A(net1029),
    .X(net1028));
 sg13g2_buf_1 fanout1029 (.A(\s0.shift_out[8] [0]),
    .X(net1029));
 sg13g2_buf_8 fanout1030 (.A(\s0.shift_out[8] [0]),
    .X(net1030));
 sg13g2_buf_8 fanout1031 (.A(net1034),
    .X(net1031));
 sg13g2_buf_8 fanout1032 (.A(net1034),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(net1034),
    .X(net1033));
 sg13g2_buf_8 fanout1034 (.A(\s0.valid_out[8] [0]),
    .X(net1034));
 sg13g2_buf_8 fanout1035 (.A(net1036),
    .X(net1035));
 sg13g2_buf_8 fanout1036 (.A(net1037),
    .X(net1036));
 sg13g2_buf_8 fanout1037 (.A(net343),
    .X(net1037));
 sg13g2_buf_8 fanout1038 (.A(net1040),
    .X(net1038));
 sg13g2_buf_1 fanout1039 (.A(net1040),
    .X(net1039));
 sg13g2_buf_8 fanout1040 (.A(\s0.shift_out[9] [0]),
    .X(net1040));
 sg13g2_buf_8 fanout1041 (.A(net1044),
    .X(net1041));
 sg13g2_buf_1 fanout1042 (.A(net1044),
    .X(net1042));
 sg13g2_buf_8 fanout1043 (.A(net1044),
    .X(net1043));
 sg13g2_buf_2 fanout1044 (.A(\s0.valid_out[9] [0]),
    .X(net1044));
 sg13g2_buf_8 fanout1045 (.A(net1048),
    .X(net1045));
 sg13g2_buf_8 fanout1046 (.A(net1048),
    .X(net1046));
 sg13g2_buf_8 fanout1047 (.A(net1048),
    .X(net1047));
 sg13g2_buf_8 fanout1048 (.A(net593),
    .X(net1048));
 sg13g2_buf_8 fanout1049 (.A(net1052),
    .X(net1049));
 sg13g2_buf_8 fanout1050 (.A(net1052),
    .X(net1050));
 sg13g2_buf_8 fanout1051 (.A(net1052),
    .X(net1051));
 sg13g2_buf_8 fanout1052 (.A(net603),
    .X(net1052));
 sg13g2_buf_8 fanout1053 (.A(net1056),
    .X(net1053));
 sg13g2_buf_2 fanout1054 (.A(net1056),
    .X(net1054));
 sg13g2_buf_8 fanout1055 (.A(net1056),
    .X(net1055));
 sg13g2_buf_8 fanout1056 (.A(net607),
    .X(net1056));
 sg13g2_buf_8 fanout1057 (.A(net1060),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(net1060),
    .X(net1058));
 sg13g2_buf_8 fanout1059 (.A(net1060),
    .X(net1059));
 sg13g2_buf_8 fanout1060 (.A(net602),
    .X(net1060));
 sg13g2_buf_8 fanout1061 (.A(net1064),
    .X(net1061));
 sg13g2_buf_8 fanout1062 (.A(net1064),
    .X(net1062));
 sg13g2_buf_8 fanout1063 (.A(net1064),
    .X(net1063));
 sg13g2_buf_8 fanout1064 (.A(net604),
    .X(net1064));
 sg13g2_buf_8 fanout1065 (.A(net1068),
    .X(net1065));
 sg13g2_buf_8 fanout1066 (.A(net1068),
    .X(net1066));
 sg13g2_buf_1 fanout1067 (.A(net1068),
    .X(net1067));
 sg13g2_buf_8 fanout1068 (.A(net600),
    .X(net1068));
 sg13g2_buf_8 fanout1069 (.A(net1072),
    .X(net1069));
 sg13g2_buf_8 fanout1070 (.A(net1072),
    .X(net1070));
 sg13g2_buf_1 fanout1071 (.A(net1072),
    .X(net1071));
 sg13g2_buf_8 fanout1072 (.A(net605),
    .X(net1072));
 sg13g2_buf_8 fanout1073 (.A(net1076),
    .X(net1073));
 sg13g2_buf_8 fanout1074 (.A(net1076),
    .X(net1074));
 sg13g2_buf_2 fanout1075 (.A(net1076),
    .X(net1075));
 sg13g2_buf_8 fanout1076 (.A(net606),
    .X(net1076));
 sg13g2_buf_8 fanout1077 (.A(net1078),
    .X(net1077));
 sg13g2_buf_8 fanout1078 (.A(net1079),
    .X(net1078));
 sg13g2_buf_8 fanout1079 (.A(net358),
    .X(net1079));
 sg13g2_buf_8 fanout1080 (.A(net1081),
    .X(net1080));
 sg13g2_buf_8 fanout1081 (.A(net1083),
    .X(net1081));
 sg13g2_buf_8 fanout1082 (.A(net1083),
    .X(net1082));
 sg13g2_buf_8 fanout1083 (.A(net358),
    .X(net1083));
 sg13g2_buf_8 fanout1084 (.A(net1087),
    .X(net1084));
 sg13g2_buf_8 fanout1085 (.A(net1087),
    .X(net1085));
 sg13g2_buf_1 fanout1086 (.A(net1087),
    .X(net1086));
 sg13g2_buf_8 fanout1087 (.A(\s0.valid_out[10] [0]),
    .X(net1087));
 sg13g2_buf_8 fanout1088 (.A(net1090),
    .X(net1088));
 sg13g2_buf_1 fanout1089 (.A(net1090),
    .X(net1089));
 sg13g2_buf_8 fanout1090 (.A(net1095),
    .X(net1090));
 sg13g2_buf_2 fanout1091 (.A(net1092),
    .X(net1091));
 sg13g2_buf_2 fanout1092 (.A(net1094),
    .X(net1092));
 sg13g2_buf_8 fanout1093 (.A(net1094),
    .X(net1093));
 sg13g2_buf_2 fanout1094 (.A(net1095),
    .X(net1094));
 sg13g2_buf_1 fanout1095 (.A(\s0.shift_out[11] [0]),
    .X(net1095));
 sg13g2_buf_8 fanout1096 (.A(net1099),
    .X(net1096));
 sg13g2_buf_8 fanout1097 (.A(net1098),
    .X(net1097));
 sg13g2_buf_8 fanout1098 (.A(net1099),
    .X(net1098));
 sg13g2_buf_8 fanout1099 (.A(net500),
    .X(net1099));
 sg13g2_buf_8 fanout1100 (.A(net1104),
    .X(net1100));
 sg13g2_buf_1 fanout1101 (.A(net1104),
    .X(net1101));
 sg13g2_buf_8 fanout1102 (.A(net1104),
    .X(net1102));
 sg13g2_buf_1 fanout1103 (.A(net1104),
    .X(net1103));
 sg13g2_buf_2 fanout1104 (.A(\s0.shift_out[12] [0]),
    .X(net1104));
 sg13g2_buf_8 fanout1105 (.A(net1106),
    .X(net1105));
 sg13g2_buf_2 fanout1106 (.A(net1107),
    .X(net1106));
 sg13g2_buf_8 fanout1107 (.A(\s0.shift_out[12] [0]),
    .X(net1107));
 sg13g2_buf_8 fanout1108 (.A(\s0.valid_out[12] [0]),
    .X(net1108));
 sg13g2_buf_1 fanout1109 (.A(\s0.valid_out[12] [0]),
    .X(net1109));
 sg13g2_buf_8 fanout1110 (.A(net1111),
    .X(net1110));
 sg13g2_buf_8 fanout1111 (.A(\s0.valid_out[12] [0]),
    .X(net1111));
 sg13g2_buf_2 fanout1112 (.A(net1113),
    .X(net1112));
 sg13g2_buf_8 fanout1113 (.A(net1116),
    .X(net1113));
 sg13g2_buf_8 fanout1114 (.A(net1116),
    .X(net1114));
 sg13g2_buf_1 fanout1115 (.A(net1116),
    .X(net1115));
 sg13g2_buf_8 fanout1116 (.A(net1118),
    .X(net1116));
 sg13g2_buf_8 fanout1117 (.A(net1118),
    .X(net1117));
 sg13g2_buf_8 fanout1118 (.A(\s0.shift_out[13] [0]),
    .X(net1118));
 sg13g2_buf_8 fanout1119 (.A(net1120),
    .X(net1119));
 sg13g2_buf_8 fanout1120 (.A(\s0.valid_out[13] [0]),
    .X(net1120));
 sg13g2_buf_8 fanout1121 (.A(\s0.valid_out[13] [0]),
    .X(net1121));
 sg13g2_buf_2 fanout1122 (.A(net1123),
    .X(net1122));
 sg13g2_buf_1 fanout1123 (.A(net1124),
    .X(net1123));
 sg13g2_buf_1 fanout1124 (.A(net1129),
    .X(net1124));
 sg13g2_buf_8 fanout1125 (.A(net1129),
    .X(net1125));
 sg13g2_buf_1 fanout1126 (.A(net1129),
    .X(net1126));
 sg13g2_buf_8 fanout1127 (.A(net1128),
    .X(net1127));
 sg13g2_buf_8 fanout1128 (.A(net1129),
    .X(net1128));
 sg13g2_buf_8 fanout1129 (.A(net335),
    .X(net1129));
 sg13g2_buf_8 fanout1130 (.A(net1133),
    .X(net1130));
 sg13g2_buf_8 fanout1131 (.A(net1133),
    .X(net1131));
 sg13g2_buf_2 fanout1132 (.A(net1133),
    .X(net1132));
 sg13g2_buf_8 fanout1133 (.A(\s0.valid_out[14] [0]),
    .X(net1133));
 sg13g2_buf_8 fanout1134 (.A(net1135),
    .X(net1134));
 sg13g2_buf_8 fanout1135 (.A(net1140),
    .X(net1135));
 sg13g2_buf_8 fanout1136 (.A(net1137),
    .X(net1136));
 sg13g2_buf_1 fanout1137 (.A(net1140),
    .X(net1137));
 sg13g2_buf_8 fanout1138 (.A(net1139),
    .X(net1138));
 sg13g2_buf_8 fanout1139 (.A(net1140),
    .X(net1139));
 sg13g2_buf_8 fanout1140 (.A(net336),
    .X(net1140));
 sg13g2_buf_8 fanout1141 (.A(net1143),
    .X(net1141));
 sg13g2_buf_8 fanout1142 (.A(net1143),
    .X(net1142));
 sg13g2_buf_8 fanout1143 (.A(net601),
    .X(net1143));
 sg13g2_buf_2 fanout1144 (.A(net1145),
    .X(net1144));
 sg13g2_buf_1 fanout1145 (.A(net1147),
    .X(net1145));
 sg13g2_buf_8 fanout1146 (.A(net1147),
    .X(net1146));
 sg13g2_buf_8 fanout1147 (.A(net1150),
    .X(net1147));
 sg13g2_buf_8 fanout1148 (.A(net1150),
    .X(net1148));
 sg13g2_buf_8 fanout1149 (.A(net1150),
    .X(net1149));
 sg13g2_buf_2 fanout1150 (.A(net338),
    .X(net1150));
 sg13g2_buf_8 fanout1151 (.A(net1154),
    .X(net1151));
 sg13g2_buf_8 fanout1152 (.A(net1154),
    .X(net1152));
 sg13g2_buf_2 fanout1153 (.A(net1154),
    .X(net1153));
 sg13g2_buf_8 fanout1154 (.A(\s0.valid_out[16] [0]),
    .X(net1154));
 sg13g2_buf_8 fanout1155 (.A(net1157),
    .X(net1155));
 sg13g2_buf_1 fanout1156 (.A(net1157),
    .X(net1156));
 sg13g2_buf_2 fanout1157 (.A(net1162),
    .X(net1157));
 sg13g2_buf_8 fanout1158 (.A(net1159),
    .X(net1158));
 sg13g2_buf_1 fanout1159 (.A(net1162),
    .X(net1159));
 sg13g2_buf_8 fanout1160 (.A(net1161),
    .X(net1160));
 sg13g2_buf_8 fanout1161 (.A(net1162),
    .X(net1161));
 sg13g2_buf_8 fanout1162 (.A(\s0.shift_out[17] [0]),
    .X(net1162));
 sg13g2_buf_8 fanout1163 (.A(net1166),
    .X(net1163));
 sg13g2_buf_8 fanout1164 (.A(net1166),
    .X(net1164));
 sg13g2_buf_2 fanout1165 (.A(net1166),
    .X(net1165));
 sg13g2_buf_8 fanout1166 (.A(\s0.valid_out[17] [0]),
    .X(net1166));
 sg13g2_buf_2 fanout1167 (.A(net1168),
    .X(net1167));
 sg13g2_buf_2 fanout1168 (.A(net1173),
    .X(net1168));
 sg13g2_buf_8 fanout1169 (.A(net1173),
    .X(net1169));
 sg13g2_buf_8 fanout1170 (.A(net1172),
    .X(net1170));
 sg13g2_buf_8 fanout1171 (.A(net1172),
    .X(net1171));
 sg13g2_buf_8 fanout1172 (.A(net1173),
    .X(net1172));
 sg13g2_buf_8 fanout1173 (.A(\s0.shift_out[18] [0]),
    .X(net1173));
 sg13g2_buf_8 fanout1174 (.A(net1177),
    .X(net1174));
 sg13g2_buf_1 fanout1175 (.A(net1177),
    .X(net1175));
 sg13g2_buf_8 fanout1176 (.A(net1177),
    .X(net1176));
 sg13g2_buf_8 fanout1177 (.A(\s0.valid_out[18] [0]),
    .X(net1177));
 sg13g2_buf_2 fanout1178 (.A(net1179),
    .X(net1178));
 sg13g2_buf_1 fanout1179 (.A(net1180),
    .X(net1179));
 sg13g2_buf_1 fanout1180 (.A(net1181),
    .X(net1180));
 sg13g2_buf_8 fanout1181 (.A(net1185),
    .X(net1181));
 sg13g2_buf_8 fanout1182 (.A(net1183),
    .X(net1182));
 sg13g2_buf_8 fanout1183 (.A(net1185),
    .X(net1183));
 sg13g2_buf_1 fanout1184 (.A(net1185),
    .X(net1184));
 sg13g2_buf_2 fanout1185 (.A(\s0.shift_out[19] [0]),
    .X(net1185));
 sg13g2_buf_8 fanout1186 (.A(net1189),
    .X(net1186));
 sg13g2_buf_1 fanout1187 (.A(net1189),
    .X(net1187));
 sg13g2_buf_8 fanout1188 (.A(net1189),
    .X(net1188));
 sg13g2_buf_8 fanout1189 (.A(net337),
    .X(net1189));
 sg13g2_buf_8 fanout1190 (.A(net1191),
    .X(net1190));
 sg13g2_buf_1 fanout1191 (.A(net1192),
    .X(net1191));
 sg13g2_buf_1 fanout1192 (.A(net1194),
    .X(net1192));
 sg13g2_buf_8 fanout1193 (.A(net1194),
    .X(net1193));
 sg13g2_buf_2 fanout1194 (.A(net333),
    .X(net1194));
 sg13g2_buf_8 fanout1195 (.A(net1196),
    .X(net1195));
 sg13g2_buf_8 fanout1196 (.A(net333),
    .X(net1196));
 sg13g2_buf_1 fanout1197 (.A(net333),
    .X(net1197));
 sg13g2_buf_8 fanout1198 (.A(net1201),
    .X(net1198));
 sg13g2_buf_1 fanout1199 (.A(net1201),
    .X(net1199));
 sg13g2_buf_8 fanout1200 (.A(net1201),
    .X(net1200));
 sg13g2_buf_2 fanout1201 (.A(\s0.valid_out[20] [0]),
    .X(net1201));
 sg13g2_buf_8 fanout1202 (.A(net1203),
    .X(net1202));
 sg13g2_buf_8 fanout1203 (.A(net332),
    .X(net1203));
 sg13g2_buf_8 fanout1204 (.A(net332),
    .X(net1204));
 sg13g2_buf_1 fanout1205 (.A(net332),
    .X(net1205));
 sg13g2_buf_8 fanout1206 (.A(net1207),
    .X(net1206));
 sg13g2_buf_8 fanout1207 (.A(\s0.valid_out[21] [0]),
    .X(net1207));
 sg13g2_buf_8 fanout1208 (.A(net1210),
    .X(net1208));
 sg13g2_buf_8 fanout1209 (.A(net1210),
    .X(net1209));
 sg13g2_buf_8 fanout1210 (.A(_2621_),
    .X(net1210));
 sg13g2_buf_8 fanout1211 (.A(net1212),
    .X(net1211));
 sg13g2_buf_8 fanout1212 (.A(_2480_),
    .X(net1212));
 sg13g2_buf_8 fanout1213 (.A(_2480_),
    .X(net1213));
 sg13g2_buf_8 fanout1214 (.A(net1215),
    .X(net1214));
 sg13g2_buf_8 fanout1215 (.A(_2476_),
    .X(net1215));
 sg13g2_buf_8 fanout1216 (.A(net1218),
    .X(net1216));
 sg13g2_buf_2 fanout1217 (.A(net1218),
    .X(net1217));
 sg13g2_buf_8 fanout1218 (.A(net1219),
    .X(net1218));
 sg13g2_buf_8 fanout1219 (.A(_2450_),
    .X(net1219));
 sg13g2_buf_8 fanout1220 (.A(_2450_),
    .X(net1220));
 sg13g2_buf_8 fanout1221 (.A(_2450_),
    .X(net1221));
 sg13g2_buf_8 fanout1222 (.A(_2449_),
    .X(net1222));
 sg13g2_buf_8 fanout1223 (.A(uio_in[1]),
    .X(net1223));
 sg13g2_buf_1 fanout1224 (.A(uio_in[1]),
    .X(net1224));
 sg13g2_buf_8 fanout1225 (.A(net1227),
    .X(net1225));
 sg13g2_buf_8 fanout1226 (.A(net1227),
    .X(net1226));
 sg13g2_buf_8 fanout1227 (.A(uio_in[0]),
    .X(net1227));
 sg13g2_buf_8 fanout1228 (.A(net1230),
    .X(net1228));
 sg13g2_buf_8 fanout1229 (.A(net1230),
    .X(net1229));
 sg13g2_buf_8 fanout1230 (.A(uio_in[0]),
    .X(net1230));
 sg13g2_buf_8 fanout1231 (.A(net1234),
    .X(net1231));
 sg13g2_buf_2 fanout1232 (.A(net1234),
    .X(net1232));
 sg13g2_buf_8 fanout1233 (.A(net1234),
    .X(net1233));
 sg13g2_buf_8 fanout1234 (.A(ui_in[7]),
    .X(net1234));
 sg13g2_buf_8 fanout1235 (.A(net1238),
    .X(net1235));
 sg13g2_buf_8 fanout1236 (.A(net1238),
    .X(net1236));
 sg13g2_buf_8 fanout1237 (.A(net1238),
    .X(net1237));
 sg13g2_buf_8 fanout1238 (.A(ui_in[7]),
    .X(net1238));
 sg13g2_buf_8 fanout1239 (.A(net1241),
    .X(net1239));
 sg13g2_buf_8 fanout1240 (.A(net1241),
    .X(net1240));
 sg13g2_buf_8 fanout1241 (.A(net1245),
    .X(net1241));
 sg13g2_buf_8 fanout1242 (.A(net1245),
    .X(net1242));
 sg13g2_buf_8 fanout1243 (.A(net1245),
    .X(net1243));
 sg13g2_buf_8 fanout1244 (.A(net1245),
    .X(net1244));
 sg13g2_buf_8 fanout1245 (.A(ui_in[6]),
    .X(net1245));
 sg13g2_buf_8 fanout1246 (.A(net1249),
    .X(net1246));
 sg13g2_buf_1 fanout1247 (.A(net1249),
    .X(net1247));
 sg13g2_buf_8 fanout1248 (.A(net1249),
    .X(net1248));
 sg13g2_buf_8 fanout1249 (.A(ui_in[5]),
    .X(net1249));
 sg13g2_buf_8 fanout1250 (.A(net1253),
    .X(net1250));
 sg13g2_buf_8 fanout1251 (.A(net1253),
    .X(net1251));
 sg13g2_buf_8 fanout1252 (.A(net1253),
    .X(net1252));
 sg13g2_buf_8 fanout1253 (.A(ui_in[5]),
    .X(net1253));
 sg13g2_buf_8 fanout1254 (.A(net1259),
    .X(net1254));
 sg13g2_buf_1 fanout1255 (.A(net1259),
    .X(net1255));
 sg13g2_buf_8 fanout1256 (.A(net1259),
    .X(net1256));
 sg13g2_buf_1 fanout1257 (.A(net1259),
    .X(net1257));
 sg13g2_buf_8 fanout1258 (.A(net1259),
    .X(net1258));
 sg13g2_buf_8 fanout1259 (.A(ui_in[4]),
    .X(net1259));
 sg13g2_buf_8 fanout1260 (.A(net1263),
    .X(net1260));
 sg13g2_buf_1 fanout1261 (.A(net1263),
    .X(net1261));
 sg13g2_buf_8 fanout1262 (.A(net1263),
    .X(net1262));
 sg13g2_buf_8 fanout1263 (.A(ui_in[3]),
    .X(net1263));
 sg13g2_buf_8 fanout1264 (.A(net1267),
    .X(net1264));
 sg13g2_buf_8 fanout1265 (.A(net1267),
    .X(net1265));
 sg13g2_buf_8 fanout1266 (.A(net1267),
    .X(net1266));
 sg13g2_buf_8 fanout1267 (.A(ui_in[3]),
    .X(net1267));
 sg13g2_buf_8 fanout1268 (.A(net1272),
    .X(net1268));
 sg13g2_buf_1 fanout1269 (.A(net1272),
    .X(net1269));
 sg13g2_buf_8 fanout1270 (.A(net1271),
    .X(net1270));
 sg13g2_buf_8 fanout1271 (.A(net1272),
    .X(net1271));
 sg13g2_buf_8 fanout1272 (.A(ui_in[2]),
    .X(net1272));
 sg13g2_buf_8 fanout1273 (.A(net1276),
    .X(net1273));
 sg13g2_buf_1 fanout1274 (.A(net1276),
    .X(net1274));
 sg13g2_buf_8 fanout1275 (.A(net1276),
    .X(net1275));
 sg13g2_buf_8 fanout1276 (.A(ui_in[1]),
    .X(net1276));
 sg13g2_buf_8 fanout1277 (.A(net1280),
    .X(net1277));
 sg13g2_buf_8 fanout1278 (.A(net1279),
    .X(net1278));
 sg13g2_buf_8 fanout1279 (.A(net1280),
    .X(net1279));
 sg13g2_buf_8 fanout1280 (.A(ui_in[1]),
    .X(net1280));
 sg13g2_buf_8 fanout1281 (.A(net1284),
    .X(net1281));
 sg13g2_buf_8 fanout1282 (.A(net1284),
    .X(net1282));
 sg13g2_buf_8 fanout1283 (.A(net1284),
    .X(net1283));
 sg13g2_buf_8 fanout1284 (.A(ui_in[0]),
    .X(net1284));
 sg13g2_buf_8 fanout1285 (.A(net1291),
    .X(net1285));
 sg13g2_buf_8 fanout1286 (.A(net1288),
    .X(net1286));
 sg13g2_buf_8 fanout1287 (.A(net1288),
    .X(net1287));
 sg13g2_buf_8 fanout1288 (.A(net1290),
    .X(net1288));
 sg13g2_buf_8 fanout1289 (.A(net1290),
    .X(net1289));
 sg13g2_buf_8 fanout1290 (.A(net1291),
    .X(net1290));
 sg13g2_buf_8 fanout1291 (.A(net1350),
    .X(net1291));
 sg13g2_buf_8 fanout1292 (.A(net1296),
    .X(net1292));
 sg13g2_buf_8 fanout1293 (.A(net1296),
    .X(net1293));
 sg13g2_buf_8 fanout1294 (.A(net1296),
    .X(net1294));
 sg13g2_buf_1 fanout1295 (.A(net1296),
    .X(net1295));
 sg13g2_buf_8 fanout1296 (.A(net1300),
    .X(net1296));
 sg13g2_buf_8 fanout1297 (.A(net1300),
    .X(net1297));
 sg13g2_buf_8 fanout1298 (.A(net1299),
    .X(net1298));
 sg13g2_buf_8 fanout1299 (.A(net1300),
    .X(net1299));
 sg13g2_buf_8 fanout1300 (.A(net1350),
    .X(net1300));
 sg13g2_buf_8 fanout1301 (.A(net1302),
    .X(net1301));
 sg13g2_buf_2 fanout1302 (.A(net1303),
    .X(net1302));
 sg13g2_buf_8 fanout1303 (.A(net1316),
    .X(net1303));
 sg13g2_buf_8 fanout1304 (.A(net1305),
    .X(net1304));
 sg13g2_buf_8 fanout1305 (.A(net1306),
    .X(net1305));
 sg13g2_buf_8 fanout1306 (.A(net1316),
    .X(net1306));
 sg13g2_buf_8 fanout1307 (.A(net1310),
    .X(net1307));
 sg13g2_buf_1 fanout1308 (.A(net1310),
    .X(net1308));
 sg13g2_buf_8 fanout1309 (.A(net1310),
    .X(net1309));
 sg13g2_buf_8 fanout1310 (.A(net1316),
    .X(net1310));
 sg13g2_buf_8 fanout1311 (.A(net1312),
    .X(net1311));
 sg13g2_buf_8 fanout1312 (.A(net1315),
    .X(net1312));
 sg13g2_buf_8 fanout1313 (.A(net1315),
    .X(net1313));
 sg13g2_buf_1 fanout1314 (.A(net1315),
    .X(net1314));
 sg13g2_buf_8 fanout1315 (.A(net1316),
    .X(net1315));
 sg13g2_buf_8 fanout1316 (.A(net1350),
    .X(net1316));
 sg13g2_buf_8 fanout1317 (.A(net1318),
    .X(net1317));
 sg13g2_buf_8 fanout1318 (.A(net1319),
    .X(net1318));
 sg13g2_buf_8 fanout1319 (.A(net1323),
    .X(net1319));
 sg13g2_buf_8 fanout1320 (.A(net1322),
    .X(net1320));
 sg13g2_buf_2 fanout1321 (.A(net1322),
    .X(net1321));
 sg13g2_buf_8 fanout1322 (.A(net1323),
    .X(net1322));
 sg13g2_buf_8 fanout1323 (.A(net1349),
    .X(net1323));
 sg13g2_buf_8 fanout1324 (.A(net1326),
    .X(net1324));
 sg13g2_buf_8 fanout1325 (.A(net1326),
    .X(net1325));
 sg13g2_buf_8 fanout1326 (.A(net1349),
    .X(net1326));
 sg13g2_buf_8 fanout1327 (.A(net1331),
    .X(net1327));
 sg13g2_buf_2 fanout1328 (.A(net1331),
    .X(net1328));
 sg13g2_buf_8 fanout1329 (.A(net1331),
    .X(net1329));
 sg13g2_buf_1 fanout1330 (.A(net1331),
    .X(net1330));
 sg13g2_buf_2 fanout1331 (.A(net1349),
    .X(net1331));
 sg13g2_buf_8 fanout1332 (.A(net1333),
    .X(net1332));
 sg13g2_buf_8 fanout1333 (.A(net1339),
    .X(net1333));
 sg13g2_buf_8 fanout1334 (.A(net1335),
    .X(net1334));
 sg13g2_buf_8 fanout1335 (.A(net1339),
    .X(net1335));
 sg13g2_buf_8 fanout1336 (.A(net1337),
    .X(net1336));
 sg13g2_buf_8 fanout1337 (.A(net1339),
    .X(net1337));
 sg13g2_buf_8 fanout1338 (.A(net1339),
    .X(net1338));
 sg13g2_buf_8 fanout1339 (.A(net1349),
    .X(net1339));
 sg13g2_buf_8 fanout1340 (.A(net1341),
    .X(net1340));
 sg13g2_buf_8 fanout1341 (.A(net1348),
    .X(net1341));
 sg13g2_buf_8 fanout1342 (.A(net1348),
    .X(net1342));
 sg13g2_buf_1 fanout1343 (.A(net1348),
    .X(net1343));
 sg13g2_buf_8 fanout1344 (.A(net1347),
    .X(net1344));
 sg13g2_buf_1 fanout1345 (.A(net1347),
    .X(net1345));
 sg13g2_buf_8 fanout1346 (.A(net1347),
    .X(net1346));
 sg13g2_buf_2 fanout1347 (.A(net1348),
    .X(net1347));
 sg13g2_buf_8 fanout1348 (.A(net1349),
    .X(net1348));
 sg13g2_buf_8 fanout1349 (.A(net1350),
    .X(net1349));
 sg13g2_buf_8 fanout1350 (.A(rst_n),
    .X(net1350));
 sg13g2_buf_1 output1 (.A(net1),
    .X(uio_out[2]));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uo_out[0]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[1]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[2]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[3]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[4]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[5]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[6]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[7]));
 sg13g2_tielo heichips25_top_sorter_10 (.L_LO(net10));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_leaf_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_leaf_2_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_leaf_36_clk));
 sg13g2_inv_2 clkload5 (.A(clknet_leaf_37_clk));
 sg13g2_inv_2 clkload6 (.A(clknet_leaf_35_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_14_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_30_clk));
 sg13g2_buf_8 clkload9 (.A(clknet_leaf_31_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_25_clk));
 sg13g2_inv_8 clkload11 (.A(clknet_leaf_28_clk));
 sg13g2_inv_2 clkload12 (.A(clknet_leaf_5_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_15_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_leaf_16_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_22_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_20_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_21_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\s0.genblk1[1].modules.bubble ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold2 (.A(\s0.genblk1[13].modules.bubble ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold3 (.A(\s0.genblk1[15].modules.bubble ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold4 (.A(\s0.genblk1[2].modules.bubble ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold5 (.A(\s0.genblk1[20].modules.bubble ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold6 (.A(\s0.genblk1[12].modules.bubble ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold7 (.A(\s0.genblk1[14].modules.bubble ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold8 (.A(\s0.genblk1[18].modules.bubble ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold9 (.A(\s0.genblk1[19].modules.bubble ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold10 (.A(\s0.genblk1[21].modules.bubble ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold11 (.A(\s0.genblk1[8].modules.bubble ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold12 (.A(\s0.genblk1[17].modules.bubble ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold13 (.A(\s0.genblk1[6].modules.bubble ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold14 (.A(\s0.genblk1[16].modules.bubble ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold15 (.A(\s0.genblk1[3].modules.bubble ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold16 (.A(\s0.module0.bubble ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold17 (.A(\s0.genblk1[7].modules.bubble ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold18 (.A(\s0.genblk1[9].modules.bubble ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold19 (.A(\s0.genblk1[10].modules.bubble ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold20 (.A(\s0.genblk1[11].modules.bubble ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold21 (.A(\s0.genblk1[4].modules.bubble ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold22 (.A(\s0.genblk1[5].modules.bubble ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold23 (.A(\s0.was_valid_out[3] [0]),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0224_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold25 (.A(\s0.was_valid_out[16] [0]),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0061_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold27 (.A(\s0.was_valid_out[19] [0]),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0025_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold29 (.A(\s0.data_out[18][4] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold30 (.A(\s0.was_valid_out[7] [0]),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0176_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold32 (.A(\s0.was_valid_out[1] [0]),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0248_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold34 (.A(\s0.data_out[11][4] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold35 (.A(_1035_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold36 (.A(\s0.shift_out[21] [0]),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold37 (.A(\s0.shift_out[20] [0]),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold38 (.A(\s0.data_out[0][7] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold39 (.A(\s0.shift_out[14] [0]),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold40 (.A(\s0.shift_out[15] [0]),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold41 (.A(\s0.valid_out[19] [0]),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold42 (.A(\s0.shift_out[16] [0]),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold43 (.A(\s0.shift_out[7] [0]),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold44 (.A(net1014),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold45 (.A(\s0.data_out[17][7] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0471_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold47 (.A(\s0.shift_out[9] [0]),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold48 (.A(\s0.data_out[0][5] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold49 (.A(\s0.data_out[0][2] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold50 (.A(\s0.was_valid_out[13] [0]),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0097_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold52 (.A(\s0.data_out[0][3] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold53 (.A(\s0.data_out[2][5] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold54 (.A(\s0.data_out[8][4] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold55 (.A(\s0.data_out[0][6] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold56 (.A(\s0.data_out[5][5] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold57 (.A(\s0.was_valid_out[4] [0]),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold58 (.A(\s0.shift_out[0] [0]),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold59 (.A(\s0.data_out[3][5] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold60 (.A(\s0.data_out[21][6] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0009_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold62 (.A(\s0.shift_out[10] [0]),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold63 (.A(\s0.data_out[21][4] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0007_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold65 (.A(\s0.data_out[21][5] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0008_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold67 (.A(\s0.was_valid_out[0] [0]),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold68 (.A(\s0.data_out[21][7] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0010_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold70 (.A(\s0.data_out[21][3] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0006_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold72 (.A(\s0.data_out[21][0] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0003_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold74 (.A(\s0.data_out[21][1] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold75 (.A(_2527_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold76 (.A(\s0.was_valid_out[21] [0]),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0001_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold78 (.A(\s0.data_out[0][4] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold79 (.A(\s0.was_valid_out[17] [0]),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0049_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold81 (.A(\s0.data_out[0][0] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold82 (.A(\s0.was_valid_out[14] [0]),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold83 (.A(\s0.was_valid_out[10] [0]),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0133_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold85 (.A(\s0.was_valid_out[15] [0]),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0073_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold87 (.A(\s0.was_valid_out[5] [0]),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0200_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold89 (.A(\s0.data_out[9][5] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold90 (.A(\s0.data_out[14][3] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold91 (.A(\s0.data_out[15][3] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold92 (.A(\s0.data_out[21][2] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold93 (.A(_2534_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold94 (.A(\s0.data_out[8][0] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold95 (.A(\s0.data_out[7][0] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold96 (.A(\s0.data_out[0][1] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold97 (.A(\s0.was_valid_out[2] [0]),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold98 (.A(\s0.data_out[1][4] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold99 (.A(\s0.data_out[20][5] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold100 (.A(\s0.data_out[1][1] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold101 (.A(_2304_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold102 (.A(\s0.was_valid_out[8] [0]),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0164_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold104 (.A(\s0.data_out[9][3] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold105 (.A(\s0.data_out[17][4] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold106 (.A(\s0.data_out[5][4] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold107 (.A(\s0.data_out[4][3] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold108 (.A(\s0.data_out[10][0] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold109 (.A(\s0.data_out[9][1] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold110 (.A(\s0.was_valid_out[18] [0]),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0037_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold112 (.A(\s0.was_valid_out[12] [0]),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0109_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold114 (.A(\s0.data_out[19][0] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold115 (.A(\s0.data_out[7][4] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold116 (.A(\s0.data_out[6][0] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold117 (.A(\s0.was_valid_out[11] [0]),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold118 (.A(\s0.data_out[19][4] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold119 (.A(\s0.data_out[5][3] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold120 (.A(\s0.data_out[16][4] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold121 (.A(\s0.data_out[2][4] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold122 (.A(\s0.data_out[10][1] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold123 (.A(\s0.data_out[7][1] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold124 (.A(\s0.data_out[3][2] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold125 (.A(\s0.data_out[3][1] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold126 (.A(\s0.data_out[16][2] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold127 (.A(\s0.data_out[6][4] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold128 (.A(\s0.data_out[2][0] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold129 (.A(_2182_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold130 (.A(\s0.data_out[2][1] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold131 (.A(_2189_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold132 (.A(\s0.data_out[9][0] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold133 (.A(\s0.data_out[10][4] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold134 (.A(\s0.data_out[13][4] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold135 (.A(\s0.data_out[15][1] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold136 (.A(\s0.data_out[5][0] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold137 (.A(\s0.data_out[4][1] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold138 (.A(\s0.data_out[8][3] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold139 (.A(\s0.was_valid_out[20] [0]),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold140 (.A(\s0.data_out[10][3] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold141 (.A(\s0.data_out[3][0] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold142 (.A(\s0.data_out[15][5] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold143 (.A(\s0.data_out[13][0] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold144 (.A(\s0.data_out[4][0] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold145 (.A(\s0.data_out[3][4] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold146 (.A(\s0.data_out[9][4] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold147 (.A(\s0.data_out[4][4] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold148 (.A(_1978_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold149 (.A(\s0.data_out[15][2] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold150 (.A(\s0.data_out[2][3] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold151 (.A(_2203_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold152 (.A(\s0.data_out[1][0] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold153 (.A(_2297_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold154 (.A(\s0.data_out[16][0] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold155 (.A(\s0.data_out[9][2] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold156 (.A(\s0.data_out[11][0] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold157 (.A(\s0.was_valid_out[9] [0]),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold158 (.A(\s0.data_out[6][3] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold159 (.A(\s0.data_out[20][1] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold160 (.A(\s0.data_out[16][5] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold161 (.A(\s0.data_out[14][0] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold162 (.A(\s0.data_out[1][2] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold163 (.A(_2311_),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold164 (.A(\s0.data_out[18][0] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold165 (.A(\s0.data_out[15][0] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold166 (.A(\s0.data_out[20][0] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold167 (.A(\s0.data_out[5][1] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold168 (.A(\s0.data_out[19][1] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold169 (.A(\s0.was_valid_out[6] [0]),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0188_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold171 (.A(\s0.data_out[7][2] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold172 (.A(\s0.data_out[17][0] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold173 (.A(\s0.data_out[20][4] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold174 (.A(\s0.data_out[4][5] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold175 (.A(\s0.data_out[13][1] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold176 (.A(\s0.data_out[12][3] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold177 (.A(\s0.data_out[12][0] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold178 (.A(\s0.data_out[15][4] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold179 (.A(\s0.data_out[19][2] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold180 (.A(\s0.data_out[16][1] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold181 (.A(\s0.data_out[13][2] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold182 (.A(\s0.data_out[18][3] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold183 (.A(\s0.data_out[1][5] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold184 (.A(\s0.data_out[17][3] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold185 (.A(\s0.data_out[10][5] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold186 (.A(\s0.data_out[8][5] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold187 (.A(_1518_),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold188 (.A(\s0.data_out[6][2] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold189 (.A(_1732_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold190 (.A(\s0.data_out[11][3] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold191 (.A(\s0.data_out[8][2] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold192 (.A(\s0.data_out[2][2] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold193 (.A(_2196_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold194 (.A(\s0.data_out[20][2] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold195 (.A(\s0.data_out[2][6] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold196 (.A(_2224_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold197 (.A(\s0.data_out[18][1] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0317_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold199 (.A(\s0.data_out[1][7] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold200 (.A(\s0.data_out[17][1] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0434_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold202 (.A(\s0.data_out[18][2] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0324_),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold204 (.A(\s0.valid_out[11] [0]),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold205 (.A(\s0.data_out[12][5] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold206 (.A(_1047_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold207 (.A(\s0.data_out[7][3] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold208 (.A(\s0.data_out[12][2] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold209 (.A(_1026_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold210 (.A(\s0.data_out[10][2] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold211 (.A(\s0.data_out[13][3] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0915_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold213 (.A(\s0.data_out[3][3] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold214 (.A(_2088_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold215 (.A(\s0.data_out[4][6] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold216 (.A(_1992_),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold217 (.A(\s0.data_out[1][3] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold218 (.A(_2318_),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold219 (.A(\s0.data_out[3][7] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold220 (.A(_2116_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold221 (.A(\s0.data_out[7][7] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold222 (.A(_1649_),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold223 (.A(\s0.data_out[6][7] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold224 (.A(_1767_),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold225 (.A(\s0.data_out[10][6] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold226 (.A(_1287_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold227 (.A(\s0.data_out[20][7] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold228 (.A(_2688_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold229 (.A(\s0.data_out[14][4] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold230 (.A(\s0.data_out[8][1] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold231 (.A(\s0.data_out[11][6] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold232 (.A(\s0.data_out[12][1] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold233 (.A(_1019_),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold234 (.A(\s0.data_out[17][2] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold235 (.A(\s0.data_out[10][7] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold236 (.A(_1294_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold237 (.A(\s0.data_out[4][2] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold238 (.A(_1964_),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold239 (.A(\s0.data_out[4][7] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold240 (.A(\s0.data_out[11][1] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold241 (.A(\s0.data_out[6][1] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold242 (.A(\s0.data_out[5][6] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold243 (.A(\s0.data_out[6][5] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold244 (.A(\s0.data_out[11][7] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold245 (.A(\s0.data_out[11][5] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold246 (.A(\s0.data_out[9][6] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold247 (.A(_1406_),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold248 (.A(\s0.data_out[7][6] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold249 (.A(_1642_),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold250 (.A(\s0.data_out[16][6] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0583_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold252 (.A(\s0.data_out[14][5] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0812_),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold254 (.A(\s0.data_out[16][3] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold255 (.A(\s0.data_out[19][6] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold256 (.A(_2796_),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold257 (.A(\s0.data_out[2][7] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold258 (.A(\s0.data_out[15][7] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0706_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold260 (.A(\s0.data_out[12][4] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold261 (.A(\s0.data_out[6][6] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold262 (.A(\s0.data_out[18][6] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0352_),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold264 (.A(\s0.data_out[20][3] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold265 (.A(_2660_),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold266 (.A(\s0.data_out[15][6] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0699_),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold268 (.A(\s0.data_out[14][1] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold269 (.A(\s0.data_out[9][7] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold270 (.A(_1413_),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold271 (.A(\s0.data_out[19][3] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold272 (.A(\s0.data_out[11][2] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold273 (.A(\s0.data_out[5][7] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold274 (.A(\s0.data_out[18][5] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0345_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold276 (.A(\s0.data_out[17][6] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold277 (.A(\s0.data_out[14][2] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold278 (.A(\s0.data_out[19][7] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold279 (.A(_2803_),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold280 (.A(\s0.data_out[3][6] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold281 (.A(\s0.data_out[14][7] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0826_),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold283 (.A(\s0.data_out[18][7] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold284 (.A(_0359_),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold285 (.A(\s0.data_out[5][2] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold286 (.A(\s0.data_out[17][5] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0462_),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold288 (.A(\s0.data_out[13][7] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0943_),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold290 (.A(\s0.data_out[19][5] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold291 (.A(\s0.data_out[8][6] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold292 (.A(\s0.data_out[12][6] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold293 (.A(\s0.data_out[7][5] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold294 (.A(\s0.data_out[1][6] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold295 (.A(\s0.data_out[16][7] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold296 (.A(\s0.data_out[20][6] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold297 (.A(\s0.data_new_delayed[7] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold298 (.A(\s0.data_out[12][7] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold299 (.A(\s0.data_out[8][7] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold300 (.A(_1532_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold301 (.A(\s0.data_out[13][6] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold302 (.A(\s0.data_out[14][6] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold303 (.A(\s0.data_out[13][5] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold304 (.A(\s0.data_new_delayed[2] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold305 (.A(\s0.valid_out[15] [0]),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold306 (.A(\s0.data_new_delayed[4] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold307 (.A(\s0.data_new_delayed[6] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold308 (.A(\s0.data_new_delayed[3] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold309 (.A(\s0.data_new_delayed[1] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold310 (.A(\s0.data_new_delayed[0] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold311 (.A(\s0.data_new_delayed[5] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold312 (.A(\s0.data_out[8][2] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold313 (.A(_1377_),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold314 (.A(\s0.data_out[8][5] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold315 (.A(\s0.data_out[2][2] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold316 (.A(\s0.data_out[12][2] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold317 (.A(\s0.data_out[11][3] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold318 (.A(_1032_),
    .X(net614));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_fill_2 FILLER_0_28 ();
 sg13g2_fill_1 FILLER_0_30 ();
 sg13g2_decap_8 FILLER_0_40 ();
 sg13g2_decap_4 FILLER_0_47 ();
 sg13g2_fill_1 FILLER_0_51 ();
 sg13g2_decap_4 FILLER_0_56 ();
 sg13g2_decap_4 FILLER_0_69 ();
 sg13g2_decap_8 FILLER_0_83 ();
 sg13g2_fill_2 FILLER_0_90 ();
 sg13g2_fill_1 FILLER_0_92 ();
 sg13g2_fill_2 FILLER_0_97 ();
 sg13g2_decap_4 FILLER_0_104 ();
 sg13g2_decap_8 FILLER_0_122 ();
 sg13g2_decap_8 FILLER_0_129 ();
 sg13g2_decap_4 FILLER_0_140 ();
 sg13g2_fill_2 FILLER_0_144 ();
 sg13g2_decap_8 FILLER_0_151 ();
 sg13g2_decap_8 FILLER_0_158 ();
 sg13g2_decap_8 FILLER_0_165 ();
 sg13g2_fill_2 FILLER_0_172 ();
 sg13g2_decap_8 FILLER_0_178 ();
 sg13g2_decap_8 FILLER_0_185 ();
 sg13g2_decap_8 FILLER_0_192 ();
 sg13g2_decap_8 FILLER_0_199 ();
 sg13g2_fill_2 FILLER_0_206 ();
 sg13g2_decap_8 FILLER_0_215 ();
 sg13g2_decap_8 FILLER_0_222 ();
 sg13g2_fill_2 FILLER_0_229 ();
 sg13g2_fill_1 FILLER_0_234 ();
 sg13g2_decap_8 FILLER_0_239 ();
 sg13g2_decap_8 FILLER_0_246 ();
 sg13g2_decap_8 FILLER_0_253 ();
 sg13g2_decap_8 FILLER_0_260 ();
 sg13g2_fill_1 FILLER_0_267 ();
 sg13g2_fill_1 FILLER_0_296 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_fill_2 FILLER_0_343 ();
 sg13g2_fill_1 FILLER_0_352 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_fill_1 FILLER_0_369 ();
 sg13g2_fill_2 FILLER_0_373 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_decap_8 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_4 FILLER_0_400 ();
 sg13g2_fill_2 FILLER_0_404 ();
 sg13g2_decap_8 FILLER_0_410 ();
 sg13g2_decap_8 FILLER_0_417 ();
 sg13g2_decap_8 FILLER_0_424 ();
 sg13g2_decap_8 FILLER_0_431 ();
 sg13g2_decap_8 FILLER_0_438 ();
 sg13g2_decap_8 FILLER_0_445 ();
 sg13g2_decap_8 FILLER_0_452 ();
 sg13g2_decap_8 FILLER_0_459 ();
 sg13g2_decap_8 FILLER_0_466 ();
 sg13g2_fill_1 FILLER_0_473 ();
 sg13g2_decap_8 FILLER_0_502 ();
 sg13g2_decap_8 FILLER_0_509 ();
 sg13g2_decap_8 FILLER_0_516 ();
 sg13g2_decap_8 FILLER_0_523 ();
 sg13g2_decap_8 FILLER_0_530 ();
 sg13g2_decap_8 FILLER_0_537 ();
 sg13g2_decap_8 FILLER_0_544 ();
 sg13g2_decap_8 FILLER_0_551 ();
 sg13g2_decap_8 FILLER_0_558 ();
 sg13g2_decap_8 FILLER_0_565 ();
 sg13g2_decap_8 FILLER_0_572 ();
 sg13g2_decap_8 FILLER_0_579 ();
 sg13g2_decap_8 FILLER_0_586 ();
 sg13g2_decap_8 FILLER_0_593 ();
 sg13g2_decap_8 FILLER_0_600 ();
 sg13g2_decap_8 FILLER_0_607 ();
 sg13g2_decap_8 FILLER_0_614 ();
 sg13g2_decap_8 FILLER_0_621 ();
 sg13g2_decap_8 FILLER_0_628 ();
 sg13g2_decap_8 FILLER_0_635 ();
 sg13g2_decap_8 FILLER_0_642 ();
 sg13g2_decap_8 FILLER_0_649 ();
 sg13g2_decap_8 FILLER_0_656 ();
 sg13g2_decap_8 FILLER_0_663 ();
 sg13g2_decap_8 FILLER_0_670 ();
 sg13g2_decap_8 FILLER_0_677 ();
 sg13g2_decap_8 FILLER_0_684 ();
 sg13g2_decap_8 FILLER_0_691 ();
 sg13g2_decap_8 FILLER_0_698 ();
 sg13g2_decap_8 FILLER_0_705 ();
 sg13g2_decap_8 FILLER_0_712 ();
 sg13g2_decap_8 FILLER_0_719 ();
 sg13g2_decap_8 FILLER_0_726 ();
 sg13g2_decap_8 FILLER_0_733 ();
 sg13g2_decap_8 FILLER_0_740 ();
 sg13g2_decap_8 FILLER_0_747 ();
 sg13g2_decap_8 FILLER_0_754 ();
 sg13g2_decap_8 FILLER_0_761 ();
 sg13g2_decap_8 FILLER_0_768 ();
 sg13g2_decap_8 FILLER_0_775 ();
 sg13g2_decap_8 FILLER_0_782 ();
 sg13g2_decap_8 FILLER_0_789 ();
 sg13g2_decap_8 FILLER_0_796 ();
 sg13g2_decap_8 FILLER_0_803 ();
 sg13g2_decap_8 FILLER_0_810 ();
 sg13g2_decap_8 FILLER_0_817 ();
 sg13g2_decap_8 FILLER_0_824 ();
 sg13g2_decap_8 FILLER_0_831 ();
 sg13g2_decap_8 FILLER_0_838 ();
 sg13g2_decap_8 FILLER_0_845 ();
 sg13g2_decap_8 FILLER_0_852 ();
 sg13g2_decap_8 FILLER_0_859 ();
 sg13g2_decap_8 FILLER_0_866 ();
 sg13g2_decap_8 FILLER_0_873 ();
 sg13g2_decap_8 FILLER_0_880 ();
 sg13g2_decap_8 FILLER_0_887 ();
 sg13g2_decap_8 FILLER_0_894 ();
 sg13g2_decap_8 FILLER_0_901 ();
 sg13g2_decap_8 FILLER_0_908 ();
 sg13g2_decap_8 FILLER_0_915 ();
 sg13g2_decap_8 FILLER_0_922 ();
 sg13g2_decap_8 FILLER_0_929 ();
 sg13g2_decap_8 FILLER_0_936 ();
 sg13g2_decap_8 FILLER_0_943 ();
 sg13g2_decap_8 FILLER_0_950 ();
 sg13g2_decap_8 FILLER_0_957 ();
 sg13g2_decap_8 FILLER_0_964 ();
 sg13g2_decap_8 FILLER_0_971 ();
 sg13g2_decap_8 FILLER_0_978 ();
 sg13g2_decap_8 FILLER_0_985 ();
 sg13g2_decap_8 FILLER_0_992 ();
 sg13g2_decap_8 FILLER_0_999 ();
 sg13g2_decap_8 FILLER_0_1006 ();
 sg13g2_decap_8 FILLER_0_1013 ();
 sg13g2_decap_8 FILLER_0_1020 ();
 sg13g2_fill_2 FILLER_0_1027 ();
 sg13g2_decap_8 FILLER_1_4 ();
 sg13g2_decap_8 FILLER_1_11 ();
 sg13g2_decap_4 FILLER_1_35 ();
 sg13g2_fill_2 FILLER_1_44 ();
 sg13g2_decap_4 FILLER_1_82 ();
 sg13g2_fill_2 FILLER_1_86 ();
 sg13g2_decap_8 FILLER_1_121 ();
 sg13g2_decap_8 FILLER_1_159 ();
 sg13g2_fill_2 FILLER_1_166 ();
 sg13g2_fill_1 FILLER_1_168 ();
 sg13g2_decap_4 FILLER_1_197 ();
 sg13g2_fill_2 FILLER_1_284 ();
 sg13g2_decap_8 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_1_436 ();
 sg13g2_decap_4 FILLER_1_443 ();
 sg13g2_fill_1 FILLER_1_475 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_4 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_522 ();
 sg13g2_decap_8 FILLER_1_529 ();
 sg13g2_decap_8 FILLER_1_536 ();
 sg13g2_decap_8 FILLER_1_543 ();
 sg13g2_decap_8 FILLER_1_550 ();
 sg13g2_decap_8 FILLER_1_557 ();
 sg13g2_decap_8 FILLER_1_564 ();
 sg13g2_decap_8 FILLER_1_571 ();
 sg13g2_decap_8 FILLER_1_578 ();
 sg13g2_decap_8 FILLER_1_585 ();
 sg13g2_decap_8 FILLER_1_592 ();
 sg13g2_decap_8 FILLER_1_599 ();
 sg13g2_decap_8 FILLER_1_606 ();
 sg13g2_decap_8 FILLER_1_613 ();
 sg13g2_decap_8 FILLER_1_620 ();
 sg13g2_decap_8 FILLER_1_627 ();
 sg13g2_decap_8 FILLER_1_634 ();
 sg13g2_decap_8 FILLER_1_641 ();
 sg13g2_decap_8 FILLER_1_648 ();
 sg13g2_decap_8 FILLER_1_655 ();
 sg13g2_decap_8 FILLER_1_662 ();
 sg13g2_decap_8 FILLER_1_669 ();
 sg13g2_decap_8 FILLER_1_676 ();
 sg13g2_decap_8 FILLER_1_683 ();
 sg13g2_decap_8 FILLER_1_690 ();
 sg13g2_decap_8 FILLER_1_697 ();
 sg13g2_decap_8 FILLER_1_704 ();
 sg13g2_decap_8 FILLER_1_711 ();
 sg13g2_decap_8 FILLER_1_718 ();
 sg13g2_decap_8 FILLER_1_725 ();
 sg13g2_decap_8 FILLER_1_732 ();
 sg13g2_decap_8 FILLER_1_739 ();
 sg13g2_decap_8 FILLER_1_746 ();
 sg13g2_decap_8 FILLER_1_753 ();
 sg13g2_decap_8 FILLER_1_760 ();
 sg13g2_decap_8 FILLER_1_767 ();
 sg13g2_decap_8 FILLER_1_774 ();
 sg13g2_decap_8 FILLER_1_781 ();
 sg13g2_decap_8 FILLER_1_788 ();
 sg13g2_decap_8 FILLER_1_795 ();
 sg13g2_decap_8 FILLER_1_802 ();
 sg13g2_decap_8 FILLER_1_809 ();
 sg13g2_decap_8 FILLER_1_816 ();
 sg13g2_decap_8 FILLER_1_823 ();
 sg13g2_decap_8 FILLER_1_830 ();
 sg13g2_decap_8 FILLER_1_837 ();
 sg13g2_decap_8 FILLER_1_844 ();
 sg13g2_decap_8 FILLER_1_851 ();
 sg13g2_decap_8 FILLER_1_858 ();
 sg13g2_decap_8 FILLER_1_865 ();
 sg13g2_decap_8 FILLER_1_872 ();
 sg13g2_decap_8 FILLER_1_879 ();
 sg13g2_decap_8 FILLER_1_886 ();
 sg13g2_decap_8 FILLER_1_893 ();
 sg13g2_decap_8 FILLER_1_900 ();
 sg13g2_decap_8 FILLER_1_907 ();
 sg13g2_decap_8 FILLER_1_914 ();
 sg13g2_decap_8 FILLER_1_921 ();
 sg13g2_decap_8 FILLER_1_928 ();
 sg13g2_decap_8 FILLER_1_935 ();
 sg13g2_decap_8 FILLER_1_942 ();
 sg13g2_decap_8 FILLER_1_949 ();
 sg13g2_decap_8 FILLER_1_956 ();
 sg13g2_decap_8 FILLER_1_963 ();
 sg13g2_decap_8 FILLER_1_970 ();
 sg13g2_decap_8 FILLER_1_977 ();
 sg13g2_decap_8 FILLER_1_984 ();
 sg13g2_decap_8 FILLER_1_991 ();
 sg13g2_decap_8 FILLER_1_998 ();
 sg13g2_decap_8 FILLER_1_1005 ();
 sg13g2_decap_8 FILLER_1_1012 ();
 sg13g2_decap_8 FILLER_1_1019 ();
 sg13g2_fill_2 FILLER_1_1026 ();
 sg13g2_fill_1 FILLER_1_1028 ();
 sg13g2_fill_1 FILLER_2_0 ();
 sg13g2_decap_4 FILLER_2_88 ();
 sg13g2_fill_2 FILLER_2_92 ();
 sg13g2_fill_2 FILLER_2_97 ();
 sg13g2_fill_1 FILLER_2_99 ();
 sg13g2_decap_4 FILLER_2_164 ();
 sg13g2_decap_8 FILLER_2_200 ();
 sg13g2_fill_2 FILLER_2_207 ();
 sg13g2_fill_1 FILLER_2_243 ();
 sg13g2_fill_1 FILLER_2_253 ();
 sg13g2_fill_1 FILLER_2_286 ();
 sg13g2_fill_2 FILLER_2_299 ();
 sg13g2_decap_8 FILLER_2_327 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_fill_1 FILLER_2_350 ();
 sg13g2_fill_2 FILLER_2_394 ();
 sg13g2_fill_1 FILLER_2_396 ();
 sg13g2_decap_8 FILLER_2_407 ();
 sg13g2_fill_2 FILLER_2_414 ();
 sg13g2_fill_2 FILLER_2_425 ();
 sg13g2_decap_8 FILLER_2_431 ();
 sg13g2_decap_8 FILLER_2_438 ();
 sg13g2_decap_8 FILLER_2_445 ();
 sg13g2_decap_4 FILLER_2_464 ();
 sg13g2_decap_4 FILLER_2_477 ();
 sg13g2_fill_2 FILLER_2_481 ();
 sg13g2_fill_2 FILLER_2_488 ();
 sg13g2_decap_4 FILLER_2_506 ();
 sg13g2_fill_1 FILLER_2_510 ();
 sg13g2_decap_8 FILLER_2_542 ();
 sg13g2_decap_8 FILLER_2_549 ();
 sg13g2_decap_8 FILLER_2_556 ();
 sg13g2_decap_8 FILLER_2_563 ();
 sg13g2_decap_8 FILLER_2_570 ();
 sg13g2_decap_4 FILLER_2_577 ();
 sg13g2_fill_2 FILLER_2_581 ();
 sg13g2_decap_4 FILLER_2_586 ();
 sg13g2_decap_8 FILLER_2_594 ();
 sg13g2_decap_8 FILLER_2_601 ();
 sg13g2_decap_8 FILLER_2_608 ();
 sg13g2_decap_8 FILLER_2_615 ();
 sg13g2_decap_8 FILLER_2_622 ();
 sg13g2_decap_8 FILLER_2_629 ();
 sg13g2_decap_8 FILLER_2_636 ();
 sg13g2_decap_4 FILLER_2_643 ();
 sg13g2_decap_8 FILLER_2_654 ();
 sg13g2_decap_8 FILLER_2_661 ();
 sg13g2_decap_8 FILLER_2_668 ();
 sg13g2_decap_8 FILLER_2_675 ();
 sg13g2_decap_8 FILLER_2_682 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_decap_8 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_2_868 ();
 sg13g2_decap_8 FILLER_2_875 ();
 sg13g2_decap_8 FILLER_2_882 ();
 sg13g2_decap_8 FILLER_2_889 ();
 sg13g2_decap_8 FILLER_2_896 ();
 sg13g2_decap_8 FILLER_2_903 ();
 sg13g2_decap_8 FILLER_2_910 ();
 sg13g2_decap_8 FILLER_2_917 ();
 sg13g2_decap_8 FILLER_2_924 ();
 sg13g2_decap_8 FILLER_2_931 ();
 sg13g2_decap_8 FILLER_2_938 ();
 sg13g2_decap_8 FILLER_2_945 ();
 sg13g2_decap_8 FILLER_2_952 ();
 sg13g2_decap_8 FILLER_2_959 ();
 sg13g2_decap_8 FILLER_2_966 ();
 sg13g2_decap_8 FILLER_2_973 ();
 sg13g2_decap_8 FILLER_2_980 ();
 sg13g2_decap_8 FILLER_2_987 ();
 sg13g2_decap_8 FILLER_2_994 ();
 sg13g2_decap_8 FILLER_2_1001 ();
 sg13g2_decap_8 FILLER_2_1008 ();
 sg13g2_decap_8 FILLER_2_1015 ();
 sg13g2_decap_8 FILLER_2_1022 ();
 sg13g2_fill_2 FILLER_3_4 ();
 sg13g2_decap_4 FILLER_3_10 ();
 sg13g2_fill_2 FILLER_3_14 ();
 sg13g2_fill_2 FILLER_3_25 ();
 sg13g2_decap_8 FILLER_3_48 ();
 sg13g2_decap_4 FILLER_3_55 ();
 sg13g2_fill_2 FILLER_3_59 ();
 sg13g2_fill_2 FILLER_3_79 ();
 sg13g2_fill_1 FILLER_3_81 ();
 sg13g2_fill_2 FILLER_3_99 ();
 sg13g2_fill_2 FILLER_3_106 ();
 sg13g2_fill_1 FILLER_3_108 ();
 sg13g2_decap_4 FILLER_3_124 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_fill_1 FILLER_3_175 ();
 sg13g2_fill_1 FILLER_3_234 ();
 sg13g2_fill_1 FILLER_3_247 ();
 sg13g2_fill_1 FILLER_3_262 ();
 sg13g2_fill_1 FILLER_3_281 ();
 sg13g2_fill_2 FILLER_3_313 ();
 sg13g2_fill_1 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_335 ();
 sg13g2_decap_8 FILLER_3_342 ();
 sg13g2_decap_4 FILLER_3_349 ();
 sg13g2_decap_8 FILLER_3_380 ();
 sg13g2_decap_4 FILLER_3_387 ();
 sg13g2_decap_8 FILLER_3_410 ();
 sg13g2_decap_4 FILLER_3_417 ();
 sg13g2_fill_1 FILLER_3_421 ();
 sg13g2_fill_1 FILLER_3_450 ();
 sg13g2_fill_1 FILLER_3_460 ();
 sg13g2_decap_8 FILLER_3_485 ();
 sg13g2_fill_1 FILLER_3_492 ();
 sg13g2_fill_1 FILLER_3_516 ();
 sg13g2_decap_8 FILLER_3_550 ();
 sg13g2_decap_8 FILLER_3_557 ();
 sg13g2_decap_4 FILLER_3_564 ();
 sg13g2_fill_2 FILLER_3_568 ();
 sg13g2_decap_4 FILLER_3_613 ();
 sg13g2_fill_2 FILLER_3_617 ();
 sg13g2_decap_4 FILLER_3_675 ();
 sg13g2_fill_2 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_712 ();
 sg13g2_decap_8 FILLER_3_719 ();
 sg13g2_decap_8 FILLER_3_726 ();
 sg13g2_decap_8 FILLER_3_733 ();
 sg13g2_decap_8 FILLER_3_740 ();
 sg13g2_decap_8 FILLER_3_747 ();
 sg13g2_decap_8 FILLER_3_754 ();
 sg13g2_decap_8 FILLER_3_761 ();
 sg13g2_decap_8 FILLER_3_768 ();
 sg13g2_decap_8 FILLER_3_775 ();
 sg13g2_decap_8 FILLER_3_782 ();
 sg13g2_decap_8 FILLER_3_789 ();
 sg13g2_decap_8 FILLER_3_796 ();
 sg13g2_decap_8 FILLER_3_803 ();
 sg13g2_decap_8 FILLER_3_810 ();
 sg13g2_decap_8 FILLER_3_817 ();
 sg13g2_decap_8 FILLER_3_824 ();
 sg13g2_decap_8 FILLER_3_831 ();
 sg13g2_decap_8 FILLER_3_838 ();
 sg13g2_decap_8 FILLER_3_845 ();
 sg13g2_decap_8 FILLER_3_852 ();
 sg13g2_decap_8 FILLER_3_859 ();
 sg13g2_decap_8 FILLER_3_866 ();
 sg13g2_decap_8 FILLER_3_873 ();
 sg13g2_decap_8 FILLER_3_880 ();
 sg13g2_decap_8 FILLER_3_887 ();
 sg13g2_decap_8 FILLER_3_894 ();
 sg13g2_decap_8 FILLER_3_901 ();
 sg13g2_decap_8 FILLER_3_908 ();
 sg13g2_decap_8 FILLER_3_915 ();
 sg13g2_decap_8 FILLER_3_922 ();
 sg13g2_decap_8 FILLER_3_929 ();
 sg13g2_decap_8 FILLER_3_936 ();
 sg13g2_decap_8 FILLER_3_943 ();
 sg13g2_decap_8 FILLER_3_950 ();
 sg13g2_decap_8 FILLER_3_957 ();
 sg13g2_decap_8 FILLER_3_964 ();
 sg13g2_decap_8 FILLER_3_971 ();
 sg13g2_decap_8 FILLER_3_978 ();
 sg13g2_decap_8 FILLER_3_985 ();
 sg13g2_decap_8 FILLER_3_992 ();
 sg13g2_decap_8 FILLER_3_999 ();
 sg13g2_decap_8 FILLER_3_1006 ();
 sg13g2_decap_8 FILLER_3_1013 ();
 sg13g2_decap_8 FILLER_3_1020 ();
 sg13g2_fill_2 FILLER_3_1027 ();
 sg13g2_decap_4 FILLER_4_4 ();
 sg13g2_fill_1 FILLER_4_8 ();
 sg13g2_decap_8 FILLER_4_13 ();
 sg13g2_fill_2 FILLER_4_20 ();
 sg13g2_fill_1 FILLER_4_22 ();
 sg13g2_fill_2 FILLER_4_27 ();
 sg13g2_fill_1 FILLER_4_29 ();
 sg13g2_fill_1 FILLER_4_39 ();
 sg13g2_decap_4 FILLER_4_55 ();
 sg13g2_decap_8 FILLER_4_78 ();
 sg13g2_decap_4 FILLER_4_85 ();
 sg13g2_fill_2 FILLER_4_116 ();
 sg13g2_fill_2 FILLER_4_126 ();
 sg13g2_fill_1 FILLER_4_128 ();
 sg13g2_decap_8 FILLER_4_134 ();
 sg13g2_decap_4 FILLER_4_141 ();
 sg13g2_fill_2 FILLER_4_145 ();
 sg13g2_decap_8 FILLER_4_152 ();
 sg13g2_fill_1 FILLER_4_159 ();
 sg13g2_fill_2 FILLER_4_188 ();
 sg13g2_fill_1 FILLER_4_190 ();
 sg13g2_fill_2 FILLER_4_205 ();
 sg13g2_fill_2 FILLER_4_224 ();
 sg13g2_decap_4 FILLER_4_259 ();
 sg13g2_decap_4 FILLER_4_288 ();
 sg13g2_fill_2 FILLER_4_292 ();
 sg13g2_fill_2 FILLER_4_314 ();
 sg13g2_decap_8 FILLER_4_340 ();
 sg13g2_fill_1 FILLER_4_347 ();
 sg13g2_decap_4 FILLER_4_373 ();
 sg13g2_fill_1 FILLER_4_377 ();
 sg13g2_decap_8 FILLER_4_382 ();
 sg13g2_fill_2 FILLER_4_401 ();
 sg13g2_fill_2 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_431 ();
 sg13g2_decap_4 FILLER_4_438 ();
 sg13g2_fill_2 FILLER_4_465 ();
 sg13g2_fill_1 FILLER_4_467 ();
 sg13g2_fill_2 FILLER_4_483 ();
 sg13g2_fill_1 FILLER_4_485 ();
 sg13g2_fill_1 FILLER_4_516 ();
 sg13g2_fill_2 FILLER_4_560 ();
 sg13g2_fill_1 FILLER_4_562 ();
 sg13g2_decap_4 FILLER_4_592 ();
 sg13g2_fill_1 FILLER_4_596 ();
 sg13g2_decap_8 FILLER_4_606 ();
 sg13g2_decap_8 FILLER_4_613 ();
 sg13g2_decap_4 FILLER_4_620 ();
 sg13g2_fill_1 FILLER_4_631 ();
 sg13g2_fill_2 FILLER_4_637 ();
 sg13g2_fill_1 FILLER_4_639 ();
 sg13g2_fill_1 FILLER_4_649 ();
 sg13g2_fill_2 FILLER_4_655 ();
 sg13g2_fill_2 FILLER_4_671 ();
 sg13g2_fill_1 FILLER_4_673 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_fill_1 FILLER_4_686 ();
 sg13g2_fill_2 FILLER_4_697 ();
 sg13g2_fill_1 FILLER_4_699 ();
 sg13g2_decap_4 FILLER_4_719 ();
 sg13g2_fill_2 FILLER_4_723 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_4 FILLER_4_749 ();
 sg13g2_fill_1 FILLER_4_753 ();
 sg13g2_decap_8 FILLER_4_761 ();
 sg13g2_decap_8 FILLER_4_768 ();
 sg13g2_decap_4 FILLER_4_775 ();
 sg13g2_fill_2 FILLER_4_779 ();
 sg13g2_decap_8 FILLER_4_809 ();
 sg13g2_decap_8 FILLER_4_816 ();
 sg13g2_decap_8 FILLER_4_823 ();
 sg13g2_decap_8 FILLER_4_830 ();
 sg13g2_decap_8 FILLER_4_837 ();
 sg13g2_decap_8 FILLER_4_844 ();
 sg13g2_decap_8 FILLER_4_851 ();
 sg13g2_decap_8 FILLER_4_858 ();
 sg13g2_decap_8 FILLER_4_865 ();
 sg13g2_decap_8 FILLER_4_872 ();
 sg13g2_decap_8 FILLER_4_879 ();
 sg13g2_decap_8 FILLER_4_886 ();
 sg13g2_decap_8 FILLER_4_893 ();
 sg13g2_decap_8 FILLER_4_900 ();
 sg13g2_decap_8 FILLER_4_907 ();
 sg13g2_decap_8 FILLER_4_914 ();
 sg13g2_decap_8 FILLER_4_921 ();
 sg13g2_decap_8 FILLER_4_928 ();
 sg13g2_decap_8 FILLER_4_935 ();
 sg13g2_decap_8 FILLER_4_942 ();
 sg13g2_decap_8 FILLER_4_949 ();
 sg13g2_decap_8 FILLER_4_956 ();
 sg13g2_decap_8 FILLER_4_963 ();
 sg13g2_decap_8 FILLER_4_970 ();
 sg13g2_decap_8 FILLER_4_977 ();
 sg13g2_decap_8 FILLER_4_984 ();
 sg13g2_decap_8 FILLER_4_991 ();
 sg13g2_decap_8 FILLER_4_998 ();
 sg13g2_decap_8 FILLER_4_1005 ();
 sg13g2_decap_8 FILLER_4_1012 ();
 sg13g2_decap_8 FILLER_4_1019 ();
 sg13g2_fill_2 FILLER_4_1026 ();
 sg13g2_fill_1 FILLER_4_1028 ();
 sg13g2_fill_1 FILLER_5_54 ();
 sg13g2_decap_8 FILLER_5_73 ();
 sg13g2_decap_4 FILLER_5_80 ();
 sg13g2_fill_2 FILLER_5_112 ();
 sg13g2_fill_1 FILLER_5_114 ();
 sg13g2_fill_2 FILLER_5_132 ();
 sg13g2_fill_1 FILLER_5_134 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_4 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_172 ();
 sg13g2_fill_2 FILLER_5_179 ();
 sg13g2_fill_1 FILLER_5_181 ();
 sg13g2_decap_8 FILLER_5_206 ();
 sg13g2_fill_2 FILLER_5_213 ();
 sg13g2_fill_1 FILLER_5_215 ();
 sg13g2_fill_1 FILLER_5_221 ();
 sg13g2_decap_8 FILLER_5_232 ();
 sg13g2_fill_2 FILLER_5_239 ();
 sg13g2_fill_1 FILLER_5_241 ();
 sg13g2_decap_4 FILLER_5_247 ();
 sg13g2_decap_8 FILLER_5_255 ();
 sg13g2_decap_8 FILLER_5_262 ();
 sg13g2_fill_2 FILLER_5_269 ();
 sg13g2_decap_8 FILLER_5_288 ();
 sg13g2_fill_2 FILLER_5_295 ();
 sg13g2_fill_1 FILLER_5_297 ();
 sg13g2_fill_1 FILLER_5_318 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_4 FILLER_5_343 ();
 sg13g2_fill_1 FILLER_5_347 ();
 sg13g2_fill_2 FILLER_5_378 ();
 sg13g2_decap_4 FILLER_5_408 ();
 sg13g2_fill_2 FILLER_5_412 ();
 sg13g2_decap_8 FILLER_5_426 ();
 sg13g2_fill_2 FILLER_5_433 ();
 sg13g2_fill_1 FILLER_5_435 ();
 sg13g2_fill_2 FILLER_5_445 ();
 sg13g2_decap_4 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_481 ();
 sg13g2_fill_2 FILLER_5_488 ();
 sg13g2_decap_8 FILLER_5_522 ();
 sg13g2_decap_8 FILLER_5_529 ();
 sg13g2_decap_8 FILLER_5_556 ();
 sg13g2_fill_2 FILLER_5_563 ();
 sg13g2_fill_1 FILLER_5_565 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_599 ();
 sg13g2_decap_4 FILLER_5_606 ();
 sg13g2_fill_1 FILLER_5_610 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_fill_1 FILLER_5_687 ();
 sg13g2_decap_8 FILLER_5_715 ();
 sg13g2_fill_2 FILLER_5_750 ();
 sg13g2_fill_2 FILLER_5_780 ();
 sg13g2_fill_1 FILLER_5_782 ();
 sg13g2_decap_8 FILLER_5_811 ();
 sg13g2_decap_8 FILLER_5_818 ();
 sg13g2_decap_8 FILLER_5_825 ();
 sg13g2_decap_8 FILLER_5_832 ();
 sg13g2_decap_8 FILLER_5_839 ();
 sg13g2_decap_8 FILLER_5_846 ();
 sg13g2_decap_8 FILLER_5_853 ();
 sg13g2_decap_8 FILLER_5_860 ();
 sg13g2_decap_8 FILLER_5_867 ();
 sg13g2_decap_8 FILLER_5_874 ();
 sg13g2_decap_8 FILLER_5_881 ();
 sg13g2_decap_8 FILLER_5_888 ();
 sg13g2_decap_8 FILLER_5_895 ();
 sg13g2_decap_8 FILLER_5_902 ();
 sg13g2_decap_8 FILLER_5_909 ();
 sg13g2_decap_8 FILLER_5_916 ();
 sg13g2_decap_8 FILLER_5_923 ();
 sg13g2_decap_8 FILLER_5_930 ();
 sg13g2_decap_8 FILLER_5_937 ();
 sg13g2_decap_8 FILLER_5_944 ();
 sg13g2_decap_8 FILLER_5_951 ();
 sg13g2_decap_8 FILLER_5_958 ();
 sg13g2_decap_8 FILLER_5_965 ();
 sg13g2_decap_8 FILLER_5_972 ();
 sg13g2_decap_8 FILLER_5_979 ();
 sg13g2_decap_8 FILLER_5_986 ();
 sg13g2_decap_8 FILLER_5_993 ();
 sg13g2_decap_8 FILLER_5_1000 ();
 sg13g2_decap_8 FILLER_5_1007 ();
 sg13g2_decap_8 FILLER_5_1014 ();
 sg13g2_decap_8 FILLER_5_1021 ();
 sg13g2_fill_1 FILLER_5_1028 ();
 sg13g2_fill_2 FILLER_6_4 ();
 sg13g2_fill_1 FILLER_6_6 ();
 sg13g2_fill_2 FILLER_6_23 ();
 sg13g2_fill_2 FILLER_6_31 ();
 sg13g2_fill_1 FILLER_6_33 ();
 sg13g2_fill_1 FILLER_6_43 ();
 sg13g2_decap_8 FILLER_6_83 ();
 sg13g2_fill_2 FILLER_6_90 ();
 sg13g2_decap_8 FILLER_6_95 ();
 sg13g2_fill_2 FILLER_6_102 ();
 sg13g2_fill_1 FILLER_6_104 ();
 sg13g2_decap_4 FILLER_6_110 ();
 sg13g2_fill_1 FILLER_6_159 ();
 sg13g2_decap_8 FILLER_6_214 ();
 sg13g2_fill_1 FILLER_6_221 ();
 sg13g2_decap_8 FILLER_6_227 ();
 sg13g2_fill_2 FILLER_6_234 ();
 sg13g2_decap_8 FILLER_6_246 ();
 sg13g2_decap_8 FILLER_6_253 ();
 sg13g2_fill_1 FILLER_6_260 ();
 sg13g2_fill_1 FILLER_6_286 ();
 sg13g2_decap_8 FILLER_6_291 ();
 sg13g2_decap_8 FILLER_6_298 ();
 sg13g2_decap_8 FILLER_6_318 ();
 sg13g2_decap_4 FILLER_6_325 ();
 sg13g2_decap_8 FILLER_6_334 ();
 sg13g2_decap_8 FILLER_6_341 ();
 sg13g2_decap_8 FILLER_6_348 ();
 sg13g2_decap_4 FILLER_6_355 ();
 sg13g2_fill_1 FILLER_6_377 ();
 sg13g2_fill_2 FILLER_6_383 ();
 sg13g2_decap_8 FILLER_6_390 ();
 sg13g2_fill_2 FILLER_6_447 ();
 sg13g2_fill_2 FILLER_6_464 ();
 sg13g2_decap_8 FILLER_6_471 ();
 sg13g2_fill_2 FILLER_6_478 ();
 sg13g2_fill_2 FILLER_6_494 ();
 sg13g2_fill_1 FILLER_6_501 ();
 sg13g2_decap_8 FILLER_6_507 ();
 sg13g2_decap_8 FILLER_6_514 ();
 sg13g2_decap_8 FILLER_6_521 ();
 sg13g2_fill_1 FILLER_6_528 ();
 sg13g2_decap_4 FILLER_6_554 ();
 sg13g2_fill_2 FILLER_6_558 ();
 sg13g2_decap_4 FILLER_6_581 ();
 sg13g2_fill_2 FILLER_6_585 ();
 sg13g2_decap_8 FILLER_6_625 ();
 sg13g2_decap_4 FILLER_6_632 ();
 sg13g2_fill_1 FILLER_6_636 ();
 sg13g2_fill_2 FILLER_6_647 ();
 sg13g2_decap_8 FILLER_6_659 ();
 sg13g2_decap_8 FILLER_6_666 ();
 sg13g2_decap_4 FILLER_6_673 ();
 sg13g2_fill_1 FILLER_6_677 ();
 sg13g2_decap_8 FILLER_6_683 ();
 sg13g2_decap_8 FILLER_6_704 ();
 sg13g2_decap_8 FILLER_6_711 ();
 sg13g2_decap_8 FILLER_6_718 ();
 sg13g2_fill_2 FILLER_6_725 ();
 sg13g2_decap_8 FILLER_6_776 ();
 sg13g2_fill_2 FILLER_6_783 ();
 sg13g2_fill_1 FILLER_6_790 ();
 sg13g2_fill_2 FILLER_6_828 ();
 sg13g2_decap_8 FILLER_6_834 ();
 sg13g2_decap_4 FILLER_6_841 ();
 sg13g2_fill_2 FILLER_6_845 ();
 sg13g2_fill_2 FILLER_6_869 ();
 sg13g2_fill_1 FILLER_6_871 ();
 sg13g2_decap_8 FILLER_6_877 ();
 sg13g2_decap_8 FILLER_6_884 ();
 sg13g2_decap_8 FILLER_6_891 ();
 sg13g2_decap_8 FILLER_6_898 ();
 sg13g2_decap_8 FILLER_6_905 ();
 sg13g2_decap_8 FILLER_6_912 ();
 sg13g2_decap_8 FILLER_6_919 ();
 sg13g2_decap_8 FILLER_6_926 ();
 sg13g2_decap_8 FILLER_6_933 ();
 sg13g2_decap_8 FILLER_6_940 ();
 sg13g2_decap_8 FILLER_6_947 ();
 sg13g2_decap_8 FILLER_6_954 ();
 sg13g2_decap_8 FILLER_6_961 ();
 sg13g2_decap_8 FILLER_6_968 ();
 sg13g2_decap_8 FILLER_6_975 ();
 sg13g2_decap_8 FILLER_6_982 ();
 sg13g2_decap_8 FILLER_6_989 ();
 sg13g2_decap_8 FILLER_6_996 ();
 sg13g2_decap_8 FILLER_6_1003 ();
 sg13g2_decap_8 FILLER_6_1010 ();
 sg13g2_decap_8 FILLER_6_1017 ();
 sg13g2_decap_4 FILLER_6_1024 ();
 sg13g2_fill_1 FILLER_6_1028 ();
 sg13g2_fill_2 FILLER_7_27 ();
 sg13g2_fill_1 FILLER_7_29 ();
 sg13g2_fill_2 FILLER_7_40 ();
 sg13g2_decap_4 FILLER_7_54 ();
 sg13g2_fill_1 FILLER_7_58 ();
 sg13g2_fill_1 FILLER_7_68 ();
 sg13g2_decap_8 FILLER_7_82 ();
 sg13g2_decap_8 FILLER_7_89 ();
 sg13g2_decap_4 FILLER_7_96 ();
 sg13g2_fill_2 FILLER_7_114 ();
 sg13g2_fill_1 FILLER_7_116 ();
 sg13g2_decap_4 FILLER_7_128 ();
 sg13g2_fill_1 FILLER_7_154 ();
 sg13g2_fill_1 FILLER_7_171 ();
 sg13g2_fill_2 FILLER_7_195 ();
 sg13g2_fill_1 FILLER_7_197 ();
 sg13g2_decap_8 FILLER_7_208 ();
 sg13g2_decap_4 FILLER_7_215 ();
 sg13g2_fill_2 FILLER_7_219 ();
 sg13g2_fill_2 FILLER_7_242 ();
 sg13g2_fill_1 FILLER_7_244 ();
 sg13g2_decap_8 FILLER_7_258 ();
 sg13g2_decap_8 FILLER_7_265 ();
 sg13g2_fill_2 FILLER_7_301 ();
 sg13g2_fill_1 FILLER_7_303 ();
 sg13g2_fill_1 FILLER_7_314 ();
 sg13g2_decap_8 FILLER_7_320 ();
 sg13g2_decap_4 FILLER_7_327 ();
 sg13g2_fill_1 FILLER_7_331 ();
 sg13g2_decap_8 FILLER_7_345 ();
 sg13g2_decap_8 FILLER_7_352 ();
 sg13g2_decap_4 FILLER_7_359 ();
 sg13g2_fill_1 FILLER_7_363 ();
 sg13g2_decap_4 FILLER_7_379 ();
 sg13g2_fill_2 FILLER_7_389 ();
 sg13g2_fill_1 FILLER_7_409 ();
 sg13g2_decap_4 FILLER_7_430 ();
 sg13g2_decap_8 FILLER_7_447 ();
 sg13g2_fill_2 FILLER_7_454 ();
 sg13g2_decap_4 FILLER_7_472 ();
 sg13g2_fill_1 FILLER_7_476 ();
 sg13g2_fill_2 FILLER_7_490 ();
 sg13g2_fill_1 FILLER_7_492 ();
 sg13g2_decap_8 FILLER_7_517 ();
 sg13g2_decap_8 FILLER_7_524 ();
 sg13g2_fill_2 FILLER_7_531 ();
 sg13g2_fill_1 FILLER_7_533 ();
 sg13g2_fill_2 FILLER_7_544 ();
 sg13g2_fill_1 FILLER_7_554 ();
 sg13g2_decap_4 FILLER_7_560 ();
 sg13g2_fill_1 FILLER_7_564 ();
 sg13g2_fill_1 FILLER_7_594 ();
 sg13g2_fill_1 FILLER_7_600 ();
 sg13g2_decap_8 FILLER_7_618 ();
 sg13g2_decap_4 FILLER_7_625 ();
 sg13g2_fill_1 FILLER_7_634 ();
 sg13g2_decap_4 FILLER_7_649 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_4 FILLER_7_686 ();
 sg13g2_fill_1 FILLER_7_690 ();
 sg13g2_fill_2 FILLER_7_742 ();
 sg13g2_fill_1 FILLER_7_744 ();
 sg13g2_decap_8 FILLER_7_775 ();
 sg13g2_fill_2 FILLER_7_782 ();
 sg13g2_decap_4 FILLER_7_803 ();
 sg13g2_fill_1 FILLER_7_807 ();
 sg13g2_decap_8 FILLER_7_817 ();
 sg13g2_fill_1 FILLER_7_824 ();
 sg13g2_fill_1 FILLER_7_852 ();
 sg13g2_decap_8 FILLER_7_908 ();
 sg13g2_decap_8 FILLER_7_915 ();
 sg13g2_decap_8 FILLER_7_922 ();
 sg13g2_decap_8 FILLER_7_929 ();
 sg13g2_decap_8 FILLER_7_936 ();
 sg13g2_decap_8 FILLER_7_943 ();
 sg13g2_decap_8 FILLER_7_950 ();
 sg13g2_decap_8 FILLER_7_957 ();
 sg13g2_decap_8 FILLER_7_964 ();
 sg13g2_decap_8 FILLER_7_971 ();
 sg13g2_decap_8 FILLER_7_978 ();
 sg13g2_decap_8 FILLER_7_985 ();
 sg13g2_decap_8 FILLER_7_992 ();
 sg13g2_decap_8 FILLER_7_999 ();
 sg13g2_decap_8 FILLER_7_1006 ();
 sg13g2_decap_8 FILLER_7_1013 ();
 sg13g2_decap_8 FILLER_7_1020 ();
 sg13g2_fill_2 FILLER_7_1027 ();
 sg13g2_fill_1 FILLER_8_4 ();
 sg13g2_decap_8 FILLER_8_9 ();
 sg13g2_fill_1 FILLER_8_16 ();
 sg13g2_decap_4 FILLER_8_49 ();
 sg13g2_fill_2 FILLER_8_53 ();
 sg13g2_decap_8 FILLER_8_68 ();
 sg13g2_decap_4 FILLER_8_75 ();
 sg13g2_fill_1 FILLER_8_79 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_fill_1 FILLER_8_126 ();
 sg13g2_fill_2 FILLER_8_136 ();
 sg13g2_fill_1 FILLER_8_138 ();
 sg13g2_fill_2 FILLER_8_144 ();
 sg13g2_fill_1 FILLER_8_146 ();
 sg13g2_decap_8 FILLER_8_156 ();
 sg13g2_decap_4 FILLER_8_163 ();
 sg13g2_fill_2 FILLER_8_167 ();
 sg13g2_fill_2 FILLER_8_205 ();
 sg13g2_fill_1 FILLER_8_207 ();
 sg13g2_decap_8 FILLER_8_213 ();
 sg13g2_fill_2 FILLER_8_220 ();
 sg13g2_fill_1 FILLER_8_226 ();
 sg13g2_fill_2 FILLER_8_230 ();
 sg13g2_decap_8 FILLER_8_237 ();
 sg13g2_decap_8 FILLER_8_244 ();
 sg13g2_fill_2 FILLER_8_251 ();
 sg13g2_decap_8 FILLER_8_258 ();
 sg13g2_decap_4 FILLER_8_265 ();
 sg13g2_fill_1 FILLER_8_269 ();
 sg13g2_fill_2 FILLER_8_288 ();
 sg13g2_decap_4 FILLER_8_300 ();
 sg13g2_fill_1 FILLER_8_304 ();
 sg13g2_decap_4 FILLER_8_324 ();
 sg13g2_decap_4 FILLER_8_361 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_4 FILLER_8_391 ();
 sg13g2_fill_2 FILLER_8_437 ();
 sg13g2_fill_2 FILLER_8_484 ();
 sg13g2_fill_1 FILLER_8_486 ();
 sg13g2_fill_2 FILLER_8_502 ();
 sg13g2_decap_8 FILLER_8_515 ();
 sg13g2_decap_8 FILLER_8_522 ();
 sg13g2_fill_2 FILLER_8_529 ();
 sg13g2_fill_2 FILLER_8_557 ();
 sg13g2_fill_1 FILLER_8_559 ();
 sg13g2_fill_2 FILLER_8_565 ();
 sg13g2_fill_1 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_573 ();
 sg13g2_fill_1 FILLER_8_589 ();
 sg13g2_fill_2 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_612 ();
 sg13g2_decap_8 FILLER_8_619 ();
 sg13g2_decap_4 FILLER_8_626 ();
 sg13g2_fill_2 FILLER_8_684 ();
 sg13g2_decap_8 FILLER_8_746 ();
 sg13g2_fill_2 FILLER_8_753 ();
 sg13g2_fill_1 FILLER_8_755 ();
 sg13g2_decap_4 FILLER_8_775 ();
 sg13g2_fill_2 FILLER_8_779 ();
 sg13g2_fill_2 FILLER_8_791 ();
 sg13g2_fill_1 FILLER_8_793 ();
 sg13g2_fill_1 FILLER_8_816 ();
 sg13g2_fill_2 FILLER_8_848 ();
 sg13g2_decap_8 FILLER_8_886 ();
 sg13g2_decap_8 FILLER_8_893 ();
 sg13g2_decap_4 FILLER_8_900 ();
 sg13g2_fill_2 FILLER_8_904 ();
 sg13g2_decap_8 FILLER_8_915 ();
 sg13g2_decap_8 FILLER_8_922 ();
 sg13g2_decap_8 FILLER_8_929 ();
 sg13g2_decap_8 FILLER_8_936 ();
 sg13g2_decap_8 FILLER_8_943 ();
 sg13g2_decap_8 FILLER_8_950 ();
 sg13g2_decap_8 FILLER_8_957 ();
 sg13g2_decap_8 FILLER_8_964 ();
 sg13g2_decap_8 FILLER_8_971 ();
 sg13g2_decap_8 FILLER_8_978 ();
 sg13g2_decap_8 FILLER_8_985 ();
 sg13g2_decap_8 FILLER_8_992 ();
 sg13g2_decap_8 FILLER_8_999 ();
 sg13g2_decap_8 FILLER_8_1006 ();
 sg13g2_decap_8 FILLER_8_1013 ();
 sg13g2_decap_8 FILLER_8_1020 ();
 sg13g2_fill_2 FILLER_8_1027 ();
 sg13g2_decap_8 FILLER_9_8 ();
 sg13g2_fill_2 FILLER_9_15 ();
 sg13g2_fill_1 FILLER_9_17 ();
 sg13g2_fill_2 FILLER_9_31 ();
 sg13g2_fill_1 FILLER_9_33 ();
 sg13g2_fill_1 FILLER_9_38 ();
 sg13g2_decap_8 FILLER_9_43 ();
 sg13g2_decap_8 FILLER_9_59 ();
 sg13g2_decap_4 FILLER_9_70 ();
 sg13g2_fill_2 FILLER_9_102 ();
 sg13g2_fill_1 FILLER_9_104 ();
 sg13g2_decap_8 FILLER_9_136 ();
 sg13g2_decap_8 FILLER_9_143 ();
 sg13g2_decap_4 FILLER_9_150 ();
 sg13g2_fill_2 FILLER_9_199 ();
 sg13g2_decap_4 FILLER_9_218 ();
 sg13g2_decap_4 FILLER_9_239 ();
 sg13g2_fill_2 FILLER_9_243 ();
 sg13g2_decap_8 FILLER_9_304 ();
 sg13g2_fill_2 FILLER_9_311 ();
 sg13g2_fill_1 FILLER_9_334 ();
 sg13g2_fill_2 FILLER_9_342 ();
 sg13g2_fill_1 FILLER_9_366 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_fill_2 FILLER_9_396 ();
 sg13g2_fill_1 FILLER_9_398 ();
 sg13g2_fill_2 FILLER_9_403 ();
 sg13g2_decap_4 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_4 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_452 ();
 sg13g2_decap_8 FILLER_9_459 ();
 sg13g2_decap_8 FILLER_9_466 ();
 sg13g2_fill_2 FILLER_9_473 ();
 sg13g2_fill_2 FILLER_9_494 ();
 sg13g2_fill_1 FILLER_9_496 ();
 sg13g2_fill_2 FILLER_9_502 ();
 sg13g2_decap_8 FILLER_9_509 ();
 sg13g2_decap_8 FILLER_9_516 ();
 sg13g2_fill_1 FILLER_9_523 ();
 sg13g2_fill_2 FILLER_9_566 ();
 sg13g2_decap_8 FILLER_9_577 ();
 sg13g2_fill_2 FILLER_9_584 ();
 sg13g2_fill_1 FILLER_9_586 ();
 sg13g2_fill_2 FILLER_9_596 ();
 sg13g2_fill_1 FILLER_9_598 ();
 sg13g2_decap_4 FILLER_9_604 ();
 sg13g2_fill_1 FILLER_9_608 ();
 sg13g2_fill_1 FILLER_9_636 ();
 sg13g2_fill_2 FILLER_9_660 ();
 sg13g2_fill_2 FILLER_9_675 ();
 sg13g2_fill_1 FILLER_9_677 ();
 sg13g2_decap_8 FILLER_9_716 ();
 sg13g2_fill_2 FILLER_9_723 ();
 sg13g2_decap_8 FILLER_9_750 ();
 sg13g2_decap_4 FILLER_9_757 ();
 sg13g2_decap_8 FILLER_9_766 ();
 sg13g2_decap_8 FILLER_9_773 ();
 sg13g2_decap_4 FILLER_9_780 ();
 sg13g2_fill_1 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_800 ();
 sg13g2_decap_4 FILLER_9_807 ();
 sg13g2_fill_1 FILLER_9_811 ();
 sg13g2_decap_8 FILLER_9_816 ();
 sg13g2_fill_1 FILLER_9_823 ();
 sg13g2_fill_2 FILLER_9_844 ();
 sg13g2_fill_1 FILLER_9_846 ();
 sg13g2_fill_1 FILLER_9_874 ();
 sg13g2_fill_1 FILLER_9_882 ();
 sg13g2_decap_8 FILLER_9_929 ();
 sg13g2_decap_8 FILLER_9_936 ();
 sg13g2_decap_8 FILLER_9_943 ();
 sg13g2_decap_8 FILLER_9_950 ();
 sg13g2_decap_8 FILLER_9_957 ();
 sg13g2_decap_8 FILLER_9_964 ();
 sg13g2_decap_8 FILLER_9_971 ();
 sg13g2_decap_8 FILLER_9_978 ();
 sg13g2_decap_8 FILLER_9_985 ();
 sg13g2_decap_8 FILLER_9_992 ();
 sg13g2_decap_8 FILLER_9_999 ();
 sg13g2_decap_8 FILLER_9_1006 ();
 sg13g2_decap_8 FILLER_9_1013 ();
 sg13g2_decap_8 FILLER_9_1020 ();
 sg13g2_fill_2 FILLER_9_1027 ();
 sg13g2_fill_1 FILLER_10_4 ();
 sg13g2_decap_4 FILLER_10_9 ();
 sg13g2_fill_1 FILLER_10_13 ();
 sg13g2_fill_2 FILLER_10_43 ();
 sg13g2_decap_8 FILLER_10_62 ();
 sg13g2_decap_8 FILLER_10_69 ();
 sg13g2_fill_2 FILLER_10_76 ();
 sg13g2_fill_1 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_129 ();
 sg13g2_decap_8 FILLER_10_136 ();
 sg13g2_decap_4 FILLER_10_143 ();
 sg13g2_fill_2 FILLER_10_167 ();
 sg13g2_decap_4 FILLER_10_173 ();
 sg13g2_fill_2 FILLER_10_177 ();
 sg13g2_fill_1 FILLER_10_206 ();
 sg13g2_decap_8 FILLER_10_212 ();
 sg13g2_decap_4 FILLER_10_219 ();
 sg13g2_fill_2 FILLER_10_223 ();
 sg13g2_decap_4 FILLER_10_260 ();
 sg13g2_fill_2 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_302 ();
 sg13g2_fill_1 FILLER_10_322 ();
 sg13g2_fill_2 FILLER_10_332 ();
 sg13g2_fill_2 FILLER_10_347 ();
 sg13g2_fill_2 FILLER_10_353 ();
 sg13g2_fill_1 FILLER_10_355 ();
 sg13g2_fill_2 FILLER_10_369 ();
 sg13g2_fill_1 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_377 ();
 sg13g2_decap_8 FILLER_10_384 ();
 sg13g2_decap_8 FILLER_10_391 ();
 sg13g2_fill_1 FILLER_10_398 ();
 sg13g2_fill_1 FILLER_10_417 ();
 sg13g2_decap_8 FILLER_10_431 ();
 sg13g2_decap_4 FILLER_10_438 ();
 sg13g2_fill_1 FILLER_10_442 ();
 sg13g2_fill_1 FILLER_10_484 ();
 sg13g2_decap_8 FILLER_10_514 ();
 sg13g2_decap_8 FILLER_10_521 ();
 sg13g2_fill_1 FILLER_10_528 ();
 sg13g2_decap_8 FILLER_10_533 ();
 sg13g2_fill_2 FILLER_10_540 ();
 sg13g2_fill_1 FILLER_10_542 ();
 sg13g2_fill_1 FILLER_10_548 ();
 sg13g2_decap_8 FILLER_10_585 ();
 sg13g2_fill_2 FILLER_10_592 ();
 sg13g2_fill_1 FILLER_10_594 ();
 sg13g2_fill_2 FILLER_10_612 ();
 sg13g2_decap_8 FILLER_10_618 ();
 sg13g2_decap_8 FILLER_10_625 ();
 sg13g2_fill_1 FILLER_10_632 ();
 sg13g2_fill_2 FILLER_10_655 ();
 sg13g2_decap_4 FILLER_10_670 ();
 sg13g2_fill_1 FILLER_10_687 ();
 sg13g2_fill_2 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_718 ();
 sg13g2_decap_8 FILLER_10_725 ();
 sg13g2_fill_1 FILLER_10_732 ();
 sg13g2_fill_2 FILLER_10_753 ();
 sg13g2_fill_1 FILLER_10_755 ();
 sg13g2_decap_4 FILLER_10_774 ();
 sg13g2_fill_2 FILLER_10_778 ();
 sg13g2_fill_1 FILLER_10_800 ();
 sg13g2_decap_8 FILLER_10_824 ();
 sg13g2_decap_8 FILLER_10_831 ();
 sg13g2_decap_4 FILLER_10_838 ();
 sg13g2_fill_2 FILLER_10_857 ();
 sg13g2_fill_2 FILLER_10_866 ();
 sg13g2_fill_2 FILLER_10_878 ();
 sg13g2_fill_1 FILLER_10_880 ();
 sg13g2_fill_2 FILLER_10_901 ();
 sg13g2_decap_8 FILLER_10_926 ();
 sg13g2_decap_8 FILLER_10_933 ();
 sg13g2_decap_8 FILLER_10_940 ();
 sg13g2_decap_8 FILLER_10_947 ();
 sg13g2_decap_8 FILLER_10_954 ();
 sg13g2_decap_8 FILLER_10_961 ();
 sg13g2_decap_8 FILLER_10_968 ();
 sg13g2_decap_8 FILLER_10_975 ();
 sg13g2_decap_8 FILLER_10_982 ();
 sg13g2_decap_8 FILLER_10_989 ();
 sg13g2_decap_8 FILLER_10_996 ();
 sg13g2_decap_8 FILLER_10_1003 ();
 sg13g2_decap_8 FILLER_10_1010 ();
 sg13g2_decap_8 FILLER_10_1017 ();
 sg13g2_decap_4 FILLER_10_1024 ();
 sg13g2_fill_1 FILLER_10_1028 ();
 sg13g2_decap_8 FILLER_11_50 ();
 sg13g2_fill_2 FILLER_11_57 ();
 sg13g2_fill_1 FILLER_11_100 ();
 sg13g2_decap_4 FILLER_11_143 ();
 sg13g2_fill_1 FILLER_11_147 ();
 sg13g2_fill_2 FILLER_11_206 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_fill_2 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_265 ();
 sg13g2_fill_2 FILLER_11_272 ();
 sg13g2_fill_1 FILLER_11_274 ();
 sg13g2_decap_4 FILLER_11_293 ();
 sg13g2_fill_2 FILLER_11_302 ();
 sg13g2_decap_8 FILLER_11_356 ();
 sg13g2_decap_4 FILLER_11_363 ();
 sg13g2_decap_4 FILLER_11_445 ();
 sg13g2_fill_2 FILLER_11_449 ();
 sg13g2_decap_4 FILLER_11_464 ();
 sg13g2_fill_2 FILLER_11_500 ();
 sg13g2_decap_8 FILLER_11_509 ();
 sg13g2_decap_4 FILLER_11_516 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_577 ();
 sg13g2_decap_4 FILLER_11_584 ();
 sg13g2_fill_1 FILLER_11_588 ();
 sg13g2_decap_4 FILLER_11_606 ();
 sg13g2_fill_1 FILLER_11_610 ();
 sg13g2_decap_4 FILLER_11_656 ();
 sg13g2_fill_2 FILLER_11_660 ();
 sg13g2_fill_2 FILLER_11_675 ();
 sg13g2_fill_2 FILLER_11_688 ();
 sg13g2_fill_1 FILLER_11_690 ();
 sg13g2_decap_8 FILLER_11_706 ();
 sg13g2_fill_2 FILLER_11_713 ();
 sg13g2_decap_8 FILLER_11_719 ();
 sg13g2_decap_8 FILLER_11_726 ();
 sg13g2_decap_8 FILLER_11_733 ();
 sg13g2_fill_1 FILLER_11_740 ();
 sg13g2_decap_8 FILLER_11_754 ();
 sg13g2_decap_8 FILLER_11_761 ();
 sg13g2_fill_2 FILLER_11_768 ();
 sg13g2_fill_1 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_803 ();
 sg13g2_fill_2 FILLER_11_814 ();
 sg13g2_fill_2 FILLER_11_821 ();
 sg13g2_fill_2 FILLER_11_831 ();
 sg13g2_fill_1 FILLER_11_833 ();
 sg13g2_decap_4 FILLER_11_857 ();
 sg13g2_fill_2 FILLER_11_866 ();
 sg13g2_fill_1 FILLER_11_868 ();
 sg13g2_decap_8 FILLER_11_874 ();
 sg13g2_decap_4 FILLER_11_886 ();
 sg13g2_fill_2 FILLER_11_907 ();
 sg13g2_decap_8 FILLER_11_946 ();
 sg13g2_decap_8 FILLER_11_953 ();
 sg13g2_decap_8 FILLER_11_960 ();
 sg13g2_decap_8 FILLER_11_967 ();
 sg13g2_decap_8 FILLER_11_974 ();
 sg13g2_decap_8 FILLER_11_981 ();
 sg13g2_decap_8 FILLER_11_988 ();
 sg13g2_decap_8 FILLER_11_995 ();
 sg13g2_decap_8 FILLER_11_1002 ();
 sg13g2_decap_8 FILLER_11_1009 ();
 sg13g2_decap_8 FILLER_11_1016 ();
 sg13g2_decap_4 FILLER_11_1023 ();
 sg13g2_fill_2 FILLER_11_1027 ();
 sg13g2_fill_2 FILLER_12_8 ();
 sg13g2_fill_1 FILLER_12_10 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_fill_2 FILLER_12_56 ();
 sg13g2_fill_2 FILLER_12_61 ();
 sg13g2_fill_1 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_68 ();
 sg13g2_fill_2 FILLER_12_75 ();
 sg13g2_decap_8 FILLER_12_81 ();
 sg13g2_fill_2 FILLER_12_88 ();
 sg13g2_fill_1 FILLER_12_90 ();
 sg13g2_fill_1 FILLER_12_105 ();
 sg13g2_fill_2 FILLER_12_116 ();
 sg13g2_fill_1 FILLER_12_118 ();
 sg13g2_fill_2 FILLER_12_146 ();
 sg13g2_fill_1 FILLER_12_148 ();
 sg13g2_fill_1 FILLER_12_172 ();
 sg13g2_decap_4 FILLER_12_205 ();
 sg13g2_decap_8 FILLER_12_243 ();
 sg13g2_decap_4 FILLER_12_250 ();
 sg13g2_fill_2 FILLER_12_254 ();
 sg13g2_decap_8 FILLER_12_296 ();
 sg13g2_fill_2 FILLER_12_303 ();
 sg13g2_fill_1 FILLER_12_305 ();
 sg13g2_decap_8 FILLER_12_338 ();
 sg13g2_decap_8 FILLER_12_345 ();
 sg13g2_decap_8 FILLER_12_352 ();
 sg13g2_fill_1 FILLER_12_364 ();
 sg13g2_fill_2 FILLER_12_393 ();
 sg13g2_fill_1 FILLER_12_395 ();
 sg13g2_decap_4 FILLER_12_420 ();
 sg13g2_fill_1 FILLER_12_424 ();
 sg13g2_decap_8 FILLER_12_435 ();
 sg13g2_decap_4 FILLER_12_442 ();
 sg13g2_fill_1 FILLER_12_446 ();
 sg13g2_fill_2 FILLER_12_479 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_4 FILLER_12_518 ();
 sg13g2_fill_1 FILLER_12_522 ();
 sg13g2_decap_4 FILLER_12_554 ();
 sg13g2_fill_2 FILLER_12_568 ();
 sg13g2_decap_8 FILLER_12_583 ();
 sg13g2_fill_2 FILLER_12_590 ();
 sg13g2_fill_2 FILLER_12_622 ();
 sg13g2_fill_1 FILLER_12_624 ();
 sg13g2_fill_1 FILLER_12_638 ();
 sg13g2_fill_1 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_669 ();
 sg13g2_fill_2 FILLER_12_676 ();
 sg13g2_fill_1 FILLER_12_678 ();
 sg13g2_fill_2 FILLER_12_689 ();
 sg13g2_fill_1 FILLER_12_691 ();
 sg13g2_fill_2 FILLER_12_754 ();
 sg13g2_fill_2 FILLER_12_761 ();
 sg13g2_fill_1 FILLER_12_763 ();
 sg13g2_fill_2 FILLER_12_773 ();
 sg13g2_fill_2 FILLER_12_790 ();
 sg13g2_decap_8 FILLER_12_796 ();
 sg13g2_decap_4 FILLER_12_803 ();
 sg13g2_decap_4 FILLER_12_859 ();
 sg13g2_fill_1 FILLER_12_863 ();
 sg13g2_decap_8 FILLER_12_877 ();
 sg13g2_fill_1 FILLER_12_884 ();
 sg13g2_fill_1 FILLER_12_894 ();
 sg13g2_decap_8 FILLER_12_936 ();
 sg13g2_decap_8 FILLER_12_943 ();
 sg13g2_decap_8 FILLER_12_950 ();
 sg13g2_decap_8 FILLER_12_957 ();
 sg13g2_decap_8 FILLER_12_964 ();
 sg13g2_decap_8 FILLER_12_971 ();
 sg13g2_decap_8 FILLER_12_978 ();
 sg13g2_decap_8 FILLER_12_985 ();
 sg13g2_decap_8 FILLER_12_992 ();
 sg13g2_decap_8 FILLER_12_999 ();
 sg13g2_decap_8 FILLER_12_1006 ();
 sg13g2_decap_8 FILLER_12_1013 ();
 sg13g2_decap_8 FILLER_12_1020 ();
 sg13g2_fill_2 FILLER_12_1027 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_29 ();
 sg13g2_fill_1 FILLER_13_44 ();
 sg13g2_fill_1 FILLER_13_58 ();
 sg13g2_fill_2 FILLER_13_86 ();
 sg13g2_fill_1 FILLER_13_88 ();
 sg13g2_fill_2 FILLER_13_125 ();
 sg13g2_fill_1 FILLER_13_127 ();
 sg13g2_decap_8 FILLER_13_142 ();
 sg13g2_fill_1 FILLER_13_149 ();
 sg13g2_fill_2 FILLER_13_186 ();
 sg13g2_decap_8 FILLER_13_242 ();
 sg13g2_decap_4 FILLER_13_249 ();
 sg13g2_fill_1 FILLER_13_253 ();
 sg13g2_fill_2 FILLER_13_307 ();
 sg13g2_fill_1 FILLER_13_309 ();
 sg13g2_fill_2 FILLER_13_319 ();
 sg13g2_fill_1 FILLER_13_321 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_347 ();
 sg13g2_decap_8 FILLER_13_354 ();
 sg13g2_decap_4 FILLER_13_361 ();
 sg13g2_fill_2 FILLER_13_365 ();
 sg13g2_fill_2 FILLER_13_394 ();
 sg13g2_fill_2 FILLER_13_426 ();
 sg13g2_decap_8 FILLER_13_445 ();
 sg13g2_decap_4 FILLER_13_452 ();
 sg13g2_fill_2 FILLER_13_461 ();
 sg13g2_fill_2 FILLER_13_489 ();
 sg13g2_decap_8 FILLER_13_508 ();
 sg13g2_fill_1 FILLER_13_515 ();
 sg13g2_fill_2 FILLER_13_529 ();
 sg13g2_decap_4 FILLER_13_535 ();
 sg13g2_fill_1 FILLER_13_539 ();
 sg13g2_fill_1 FILLER_13_585 ();
 sg13g2_decap_4 FILLER_13_601 ();
 sg13g2_fill_2 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_643 ();
 sg13g2_decap_4 FILLER_13_650 ();
 sg13g2_fill_1 FILLER_13_654 ();
 sg13g2_decap_8 FILLER_13_674 ();
 sg13g2_fill_2 FILLER_13_681 ();
 sg13g2_fill_2 FILLER_13_692 ();
 sg13g2_decap_8 FILLER_13_719 ();
 sg13g2_decap_8 FILLER_13_726 ();
 sg13g2_decap_8 FILLER_13_733 ();
 sg13g2_fill_2 FILLER_13_740 ();
 sg13g2_fill_1 FILLER_13_780 ();
 sg13g2_fill_2 FILLER_13_829 ();
 sg13g2_fill_1 FILLER_13_831 ();
 sg13g2_fill_2 FILLER_13_860 ();
 sg13g2_decap_4 FILLER_13_881 ();
 sg13g2_fill_1 FILLER_13_912 ();
 sg13g2_decap_8 FILLER_13_917 ();
 sg13g2_decap_8 FILLER_13_928 ();
 sg13g2_decap_8 FILLER_13_935 ();
 sg13g2_decap_8 FILLER_13_942 ();
 sg13g2_decap_8 FILLER_13_949 ();
 sg13g2_decap_8 FILLER_13_956 ();
 sg13g2_decap_8 FILLER_13_963 ();
 sg13g2_decap_8 FILLER_13_970 ();
 sg13g2_decap_8 FILLER_13_977 ();
 sg13g2_decap_8 FILLER_13_984 ();
 sg13g2_decap_8 FILLER_13_991 ();
 sg13g2_decap_8 FILLER_13_998 ();
 sg13g2_decap_8 FILLER_13_1005 ();
 sg13g2_decap_8 FILLER_13_1012 ();
 sg13g2_decap_8 FILLER_13_1019 ();
 sg13g2_fill_2 FILLER_13_1026 ();
 sg13g2_fill_1 FILLER_13_1028 ();
 sg13g2_fill_2 FILLER_14_4 ();
 sg13g2_fill_2 FILLER_14_40 ();
 sg13g2_decap_8 FILLER_14_61 ();
 sg13g2_fill_2 FILLER_14_68 ();
 sg13g2_decap_4 FILLER_14_106 ();
 sg13g2_decap_4 FILLER_14_116 ();
 sg13g2_fill_2 FILLER_14_125 ();
 sg13g2_fill_2 FILLER_14_137 ();
 sg13g2_fill_2 FILLER_14_148 ();
 sg13g2_fill_2 FILLER_14_183 ();
 sg13g2_fill_1 FILLER_14_185 ();
 sg13g2_fill_1 FILLER_14_199 ();
 sg13g2_fill_1 FILLER_14_207 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_fill_2 FILLER_14_224 ();
 sg13g2_fill_1 FILLER_14_226 ();
 sg13g2_fill_2 FILLER_14_231 ();
 sg13g2_fill_1 FILLER_14_233 ();
 sg13g2_fill_2 FILLER_14_284 ();
 sg13g2_fill_1 FILLER_14_312 ();
 sg13g2_decap_4 FILLER_14_333 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_fill_2 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_fill_2 FILLER_14_413 ();
 sg13g2_fill_1 FILLER_14_415 ();
 sg13g2_decap_4 FILLER_14_429 ();
 sg13g2_fill_2 FILLER_14_433 ();
 sg13g2_decap_4 FILLER_14_479 ();
 sg13g2_fill_1 FILLER_14_483 ();
 sg13g2_fill_2 FILLER_14_494 ();
 sg13g2_decap_8 FILLER_14_501 ();
 sg13g2_fill_2 FILLER_14_508 ();
 sg13g2_fill_1 FILLER_14_510 ();
 sg13g2_decap_8 FILLER_14_515 ();
 sg13g2_fill_2 FILLER_14_522 ();
 sg13g2_fill_1 FILLER_14_524 ();
 sg13g2_fill_2 FILLER_14_552 ();
 sg13g2_fill_1 FILLER_14_554 ();
 sg13g2_decap_8 FILLER_14_565 ();
 sg13g2_fill_2 FILLER_14_572 ();
 sg13g2_decap_8 FILLER_14_579 ();
 sg13g2_fill_2 FILLER_14_586 ();
 sg13g2_fill_2 FILLER_14_598 ();
 sg13g2_decap_4 FILLER_14_627 ();
 sg13g2_fill_2 FILLER_14_651 ();
 sg13g2_fill_1 FILLER_14_653 ();
 sg13g2_fill_1 FILLER_14_667 ();
 sg13g2_decap_8 FILLER_14_678 ();
 sg13g2_decap_8 FILLER_14_685 ();
 sg13g2_fill_2 FILLER_14_727 ();
 sg13g2_fill_1 FILLER_14_729 ();
 sg13g2_decap_8 FILLER_14_734 ();
 sg13g2_decap_8 FILLER_14_741 ();
 sg13g2_fill_1 FILLER_14_752 ();
 sg13g2_decap_8 FILLER_14_758 ();
 sg13g2_decap_4 FILLER_14_765 ();
 sg13g2_fill_2 FILLER_14_769 ();
 sg13g2_fill_2 FILLER_14_781 ();
 sg13g2_fill_1 FILLER_14_783 ();
 sg13g2_fill_2 FILLER_14_797 ();
 sg13g2_decap_4 FILLER_14_832 ();
 sg13g2_fill_1 FILLER_14_836 ();
 sg13g2_decap_4 FILLER_14_841 ();
 sg13g2_fill_1 FILLER_14_852 ();
 sg13g2_fill_2 FILLER_14_862 ();
 sg13g2_fill_1 FILLER_14_864 ();
 sg13g2_fill_1 FILLER_14_873 ();
 sg13g2_decap_8 FILLER_14_884 ();
 sg13g2_decap_8 FILLER_14_901 ();
 sg13g2_decap_4 FILLER_14_908 ();
 sg13g2_fill_2 FILLER_14_912 ();
 sg13g2_fill_2 FILLER_14_923 ();
 sg13g2_fill_1 FILLER_14_925 ();
 sg13g2_decap_8 FILLER_14_954 ();
 sg13g2_decap_8 FILLER_14_961 ();
 sg13g2_decap_8 FILLER_14_968 ();
 sg13g2_decap_8 FILLER_14_975 ();
 sg13g2_decap_8 FILLER_14_982 ();
 sg13g2_decap_8 FILLER_14_989 ();
 sg13g2_decap_8 FILLER_14_996 ();
 sg13g2_decap_8 FILLER_14_1003 ();
 sg13g2_decap_8 FILLER_14_1010 ();
 sg13g2_decap_8 FILLER_14_1017 ();
 sg13g2_decap_4 FILLER_14_1024 ();
 sg13g2_fill_1 FILLER_14_1028 ();
 sg13g2_fill_1 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_42 ();
 sg13g2_fill_2 FILLER_15_48 ();
 sg13g2_fill_1 FILLER_15_50 ();
 sg13g2_decap_4 FILLER_15_56 ();
 sg13g2_fill_2 FILLER_15_65 ();
 sg13g2_fill_1 FILLER_15_67 ();
 sg13g2_fill_2 FILLER_15_93 ();
 sg13g2_fill_1 FILLER_15_95 ();
 sg13g2_decap_8 FILLER_15_134 ();
 sg13g2_decap_8 FILLER_15_146 ();
 sg13g2_fill_1 FILLER_15_198 ();
 sg13g2_decap_4 FILLER_15_211 ();
 sg13g2_fill_2 FILLER_15_225 ();
 sg13g2_fill_1 FILLER_15_227 ();
 sg13g2_decap_8 FILLER_15_232 ();
 sg13g2_decap_8 FILLER_15_246 ();
 sg13g2_decap_8 FILLER_15_253 ();
 sg13g2_decap_8 FILLER_15_260 ();
 sg13g2_decap_8 FILLER_15_267 ();
 sg13g2_decap_4 FILLER_15_274 ();
 sg13g2_fill_2 FILLER_15_291 ();
 sg13g2_decap_8 FILLER_15_303 ();
 sg13g2_fill_2 FILLER_15_310 ();
 sg13g2_fill_1 FILLER_15_312 ();
 sg13g2_fill_2 FILLER_15_327 ();
 sg13g2_fill_1 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_335 ();
 sg13g2_fill_1 FILLER_15_342 ();
 sg13g2_fill_2 FILLER_15_352 ();
 sg13g2_fill_2 FILLER_15_373 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_fill_2 FILLER_15_401 ();
 sg13g2_decap_4 FILLER_15_417 ();
 sg13g2_fill_2 FILLER_15_421 ();
 sg13g2_decap_8 FILLER_15_433 ();
 sg13g2_fill_2 FILLER_15_440 ();
 sg13g2_decap_4 FILLER_15_446 ();
 sg13g2_fill_2 FILLER_15_450 ();
 sg13g2_fill_1 FILLER_15_461 ();
 sg13g2_fill_1 FILLER_15_477 ();
 sg13g2_decap_4 FILLER_15_501 ();
 sg13g2_fill_2 FILLER_15_557 ();
 sg13g2_fill_1 FILLER_15_559 ();
 sg13g2_decap_8 FILLER_15_571 ();
 sg13g2_decap_8 FILLER_15_578 ();
 sg13g2_fill_2 FILLER_15_594 ();
 sg13g2_fill_1 FILLER_15_596 ();
 sg13g2_decap_8 FILLER_15_610 ();
 sg13g2_fill_1 FILLER_15_617 ();
 sg13g2_fill_2 FILLER_15_622 ();
 sg13g2_decap_8 FILLER_15_641 ();
 sg13g2_decap_8 FILLER_15_648 ();
 sg13g2_fill_1 FILLER_15_655 ();
 sg13g2_fill_2 FILLER_15_678 ();
 sg13g2_decap_4 FILLER_15_685 ();
 sg13g2_fill_2 FILLER_15_689 ();
 sg13g2_decap_4 FILLER_15_696 ();
 sg13g2_decap_8 FILLER_15_715 ();
 sg13g2_fill_2 FILLER_15_722 ();
 sg13g2_decap_4 FILLER_15_752 ();
 sg13g2_fill_1 FILLER_15_774 ();
 sg13g2_decap_4 FILLER_15_785 ();
 sg13g2_decap_8 FILLER_15_811 ();
 sg13g2_decap_4 FILLER_15_818 ();
 sg13g2_fill_1 FILLER_15_822 ();
 sg13g2_decap_8 FILLER_15_868 ();
 sg13g2_fill_1 FILLER_15_875 ();
 sg13g2_fill_2 FILLER_15_903 ();
 sg13g2_fill_2 FILLER_15_936 ();
 sg13g2_fill_1 FILLER_15_938 ();
 sg13g2_decap_8 FILLER_15_980 ();
 sg13g2_decap_8 FILLER_15_987 ();
 sg13g2_decap_8 FILLER_15_994 ();
 sg13g2_decap_8 FILLER_15_1001 ();
 sg13g2_decap_8 FILLER_15_1008 ();
 sg13g2_decap_8 FILLER_15_1015 ();
 sg13g2_decap_8 FILLER_15_1022 ();
 sg13g2_fill_2 FILLER_16_4 ();
 sg13g2_decap_8 FILLER_16_10 ();
 sg13g2_fill_2 FILLER_16_17 ();
 sg13g2_decap_4 FILLER_16_53 ();
 sg13g2_decap_8 FILLER_16_61 ();
 sg13g2_decap_8 FILLER_16_68 ();
 sg13g2_fill_1 FILLER_16_75 ();
 sg13g2_decap_4 FILLER_16_104 ();
 sg13g2_fill_1 FILLER_16_108 ();
 sg13g2_fill_2 FILLER_16_114 ();
 sg13g2_decap_8 FILLER_16_136 ();
 sg13g2_decap_8 FILLER_16_143 ();
 sg13g2_fill_1 FILLER_16_150 ();
 sg13g2_decap_8 FILLER_16_164 ();
 sg13g2_fill_2 FILLER_16_175 ();
 sg13g2_fill_1 FILLER_16_177 ();
 sg13g2_decap_4 FILLER_16_182 ();
 sg13g2_fill_2 FILLER_16_186 ();
 sg13g2_decap_8 FILLER_16_191 ();
 sg13g2_decap_4 FILLER_16_198 ();
 sg13g2_fill_2 FILLER_16_202 ();
 sg13g2_fill_1 FILLER_16_260 ();
 sg13g2_fill_1 FILLER_16_274 ();
 sg13g2_decap_4 FILLER_16_289 ();
 sg13g2_fill_1 FILLER_16_293 ();
 sg13g2_fill_2 FILLER_16_316 ();
 sg13g2_fill_2 FILLER_16_323 ();
 sg13g2_fill_1 FILLER_16_325 ();
 sg13g2_fill_1 FILLER_16_336 ();
 sg13g2_fill_2 FILLER_16_346 ();
 sg13g2_fill_1 FILLER_16_358 ();
 sg13g2_decap_8 FILLER_16_386 ();
 sg13g2_fill_2 FILLER_16_393 ();
 sg13g2_fill_1 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_fill_2 FILLER_16_434 ();
 sg13g2_fill_1 FILLER_16_436 ();
 sg13g2_fill_1 FILLER_16_488 ();
 sg13g2_decap_8 FILLER_16_499 ();
 sg13g2_fill_2 FILLER_16_506 ();
 sg13g2_decap_8 FILLER_16_517 ();
 sg13g2_decap_4 FILLER_16_524 ();
 sg13g2_fill_2 FILLER_16_536 ();
 sg13g2_decap_8 FILLER_16_543 ();
 sg13g2_decap_8 FILLER_16_578 ();
 sg13g2_decap_8 FILLER_16_585 ();
 sg13g2_fill_2 FILLER_16_592 ();
 sg13g2_decap_8 FILLER_16_598 ();
 sg13g2_fill_2 FILLER_16_605 ();
 sg13g2_decap_4 FILLER_16_611 ();
 sg13g2_decap_8 FILLER_16_625 ();
 sg13g2_decap_4 FILLER_16_659 ();
 sg13g2_fill_2 FILLER_16_683 ();
 sg13g2_decap_8 FILLER_16_708 ();
 sg13g2_decap_8 FILLER_16_715 ();
 sg13g2_decap_8 FILLER_16_722 ();
 sg13g2_fill_1 FILLER_16_729 ();
 sg13g2_decap_4 FILLER_16_733 ();
 sg13g2_fill_1 FILLER_16_737 ();
 sg13g2_fill_1 FILLER_16_752 ();
 sg13g2_decap_8 FILLER_16_773 ();
 sg13g2_decap_4 FILLER_16_780 ();
 sg13g2_decap_4 FILLER_16_808 ();
 sg13g2_decap_8 FILLER_16_837 ();
 sg13g2_decap_4 FILLER_16_844 ();
 sg13g2_fill_1 FILLER_16_848 ();
 sg13g2_fill_2 FILLER_16_916 ();
 sg13g2_fill_1 FILLER_16_918 ();
 sg13g2_fill_1 FILLER_16_941 ();
 sg13g2_fill_2 FILLER_16_945 ();
 sg13g2_fill_2 FILLER_16_952 ();
 sg13g2_decap_8 FILLER_16_961 ();
 sg13g2_fill_2 FILLER_16_968 ();
 sg13g2_decap_8 FILLER_16_979 ();
 sg13g2_decap_8 FILLER_16_986 ();
 sg13g2_decap_8 FILLER_16_993 ();
 sg13g2_decap_8 FILLER_16_1000 ();
 sg13g2_decap_8 FILLER_16_1007 ();
 sg13g2_decap_8 FILLER_16_1014 ();
 sg13g2_decap_8 FILLER_16_1021 ();
 sg13g2_fill_1 FILLER_16_1028 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_2 ();
 sg13g2_decap_8 FILLER_17_68 ();
 sg13g2_decap_8 FILLER_17_75 ();
 sg13g2_decap_8 FILLER_17_82 ();
 sg13g2_fill_2 FILLER_17_94 ();
 sg13g2_decap_8 FILLER_17_110 ();
 sg13g2_decap_4 FILLER_17_117 ();
 sg13g2_decap_8 FILLER_17_136 ();
 sg13g2_decap_4 FILLER_17_143 ();
 sg13g2_fill_2 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_4 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_197 ();
 sg13g2_fill_2 FILLER_17_204 ();
 sg13g2_fill_2 FILLER_17_216 ();
 sg13g2_fill_1 FILLER_17_218 ();
 sg13g2_fill_2 FILLER_17_238 ();
 sg13g2_fill_1 FILLER_17_240 ();
 sg13g2_decap_8 FILLER_17_246 ();
 sg13g2_decap_8 FILLER_17_253 ();
 sg13g2_fill_2 FILLER_17_260 ();
 sg13g2_fill_1 FILLER_17_294 ();
 sg13g2_fill_2 FILLER_17_341 ();
 sg13g2_decap_4 FILLER_17_354 ();
 sg13g2_fill_2 FILLER_17_358 ();
 sg13g2_decap_4 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_4 FILLER_17_399 ();
 sg13g2_fill_1 FILLER_17_403 ();
 sg13g2_fill_1 FILLER_17_423 ();
 sg13g2_fill_2 FILLER_17_436 ();
 sg13g2_decap_8 FILLER_17_451 ();
 sg13g2_fill_1 FILLER_17_458 ();
 sg13g2_fill_1 FILLER_17_469 ();
 sg13g2_fill_2 FILLER_17_480 ();
 sg13g2_decap_4 FILLER_17_496 ();
 sg13g2_fill_1 FILLER_17_500 ();
 sg13g2_decap_8 FILLER_17_520 ();
 sg13g2_decap_8 FILLER_17_554 ();
 sg13g2_fill_2 FILLER_17_561 ();
 sg13g2_decap_8 FILLER_17_582 ();
 sg13g2_fill_1 FILLER_17_599 ();
 sg13g2_fill_2 FILLER_17_615 ();
 sg13g2_fill_1 FILLER_17_617 ();
 sg13g2_decap_4 FILLER_17_633 ();
 sg13g2_fill_1 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_642 ();
 sg13g2_fill_1 FILLER_17_649 ();
 sg13g2_fill_2 FILLER_17_672 ();
 sg13g2_fill_2 FILLER_17_678 ();
 sg13g2_fill_1 FILLER_17_680 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_4 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_743 ();
 sg13g2_decap_8 FILLER_17_767 ();
 sg13g2_decap_4 FILLER_17_774 ();
 sg13g2_fill_1 FILLER_17_778 ();
 sg13g2_fill_2 FILLER_17_796 ();
 sg13g2_decap_8 FILLER_17_808 ();
 sg13g2_decap_8 FILLER_17_815 ();
 sg13g2_fill_2 FILLER_17_822 ();
 sg13g2_fill_1 FILLER_17_824 ();
 sg13g2_decap_8 FILLER_17_839 ();
 sg13g2_fill_1 FILLER_17_846 ();
 sg13g2_fill_2 FILLER_17_856 ();
 sg13g2_decap_8 FILLER_17_862 ();
 sg13g2_decap_8 FILLER_17_869 ();
 sg13g2_decap_4 FILLER_17_876 ();
 sg13g2_fill_2 FILLER_17_880 ();
 sg13g2_fill_2 FILLER_17_900 ();
 sg13g2_fill_1 FILLER_17_907 ();
 sg13g2_decap_8 FILLER_17_927 ();
 sg13g2_fill_1 FILLER_17_934 ();
 sg13g2_decap_8 FILLER_17_963 ();
 sg13g2_decap_8 FILLER_17_970 ();
 sg13g2_decap_8 FILLER_17_977 ();
 sg13g2_decap_8 FILLER_17_984 ();
 sg13g2_decap_8 FILLER_17_991 ();
 sg13g2_decap_8 FILLER_17_998 ();
 sg13g2_decap_8 FILLER_17_1005 ();
 sg13g2_decap_8 FILLER_17_1012 ();
 sg13g2_decap_8 FILLER_17_1019 ();
 sg13g2_fill_2 FILLER_17_1026 ();
 sg13g2_fill_1 FILLER_17_1028 ();
 sg13g2_decap_8 FILLER_18_12 ();
 sg13g2_decap_8 FILLER_18_19 ();
 sg13g2_decap_8 FILLER_18_26 ();
 sg13g2_fill_1 FILLER_18_33 ();
 sg13g2_fill_2 FILLER_18_38 ();
 sg13g2_fill_1 FILLER_18_40 ();
 sg13g2_fill_2 FILLER_18_68 ();
 sg13g2_decap_4 FILLER_18_110 ();
 sg13g2_fill_1 FILLER_18_114 ();
 sg13g2_decap_8 FILLER_18_160 ();
 sg13g2_decap_4 FILLER_18_167 ();
 sg13g2_fill_2 FILLER_18_171 ();
 sg13g2_decap_4 FILLER_18_178 ();
 sg13g2_fill_1 FILLER_18_182 ();
 sg13g2_decap_4 FILLER_18_245 ();
 sg13g2_fill_1 FILLER_18_249 ();
 sg13g2_fill_1 FILLER_18_266 ();
 sg13g2_fill_2 FILLER_18_281 ();
 sg13g2_decap_8 FILLER_18_293 ();
 sg13g2_decap_8 FILLER_18_300 ();
 sg13g2_decap_4 FILLER_18_307 ();
 sg13g2_fill_1 FILLER_18_311 ();
 sg13g2_fill_1 FILLER_18_317 ();
 sg13g2_decap_4 FILLER_18_336 ();
 sg13g2_fill_1 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_fill_2 FILLER_18_409 ();
 sg13g2_fill_1 FILLER_18_411 ();
 sg13g2_decap_8 FILLER_18_440 ();
 sg13g2_decap_4 FILLER_18_447 ();
 sg13g2_fill_1 FILLER_18_451 ();
 sg13g2_fill_2 FILLER_18_475 ();
 sg13g2_fill_2 FILLER_18_487 ();
 sg13g2_decap_8 FILLER_18_519 ();
 sg13g2_decap_8 FILLER_18_526 ();
 sg13g2_decap_8 FILLER_18_537 ();
 sg13g2_fill_2 FILLER_18_544 ();
 sg13g2_fill_1 FILLER_18_546 ();
 sg13g2_decap_8 FILLER_18_604 ();
 sg13g2_decap_4 FILLER_18_611 ();
 sg13g2_decap_8 FILLER_18_625 ();
 sg13g2_fill_2 FILLER_18_662 ();
 sg13g2_decap_8 FILLER_18_708 ();
 sg13g2_decap_4 FILLER_18_715 ();
 sg13g2_fill_1 FILLER_18_719 ();
 sg13g2_fill_1 FILLER_18_740 ();
 sg13g2_fill_1 FILLER_18_753 ();
 sg13g2_fill_1 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_781 ();
 sg13g2_fill_1 FILLER_18_798 ();
 sg13g2_fill_2 FILLER_18_813 ();
 sg13g2_fill_1 FILLER_18_815 ();
 sg13g2_fill_1 FILLER_18_848 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_18_867 ();
 sg13g2_decap_8 FILLER_18_874 ();
 sg13g2_decap_8 FILLER_18_881 ();
 sg13g2_fill_2 FILLER_18_888 ();
 sg13g2_fill_1 FILLER_18_893 ();
 sg13g2_fill_2 FILLER_18_899 ();
 sg13g2_fill_1 FILLER_18_901 ();
 sg13g2_decap_4 FILLER_18_927 ();
 sg13g2_decap_8 FILLER_18_966 ();
 sg13g2_decap_8 FILLER_18_973 ();
 sg13g2_decap_8 FILLER_18_980 ();
 sg13g2_decap_8 FILLER_18_987 ();
 sg13g2_decap_8 FILLER_18_994 ();
 sg13g2_decap_8 FILLER_18_1001 ();
 sg13g2_decap_8 FILLER_18_1008 ();
 sg13g2_decap_8 FILLER_18_1015 ();
 sg13g2_decap_8 FILLER_18_1022 ();
 sg13g2_fill_1 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_29 ();
 sg13g2_decap_8 FILLER_19_36 ();
 sg13g2_decap_8 FILLER_19_43 ();
 sg13g2_fill_2 FILLER_19_50 ();
 sg13g2_decap_4 FILLER_19_71 ();
 sg13g2_fill_1 FILLER_19_75 ();
 sg13g2_fill_2 FILLER_19_86 ();
 sg13g2_decap_8 FILLER_19_92 ();
 sg13g2_decap_8 FILLER_19_99 ();
 sg13g2_decap_8 FILLER_19_106 ();
 sg13g2_decap_4 FILLER_19_138 ();
 sg13g2_decap_4 FILLER_19_166 ();
 sg13g2_decap_8 FILLER_19_174 ();
 sg13g2_fill_2 FILLER_19_181 ();
 sg13g2_fill_1 FILLER_19_183 ();
 sg13g2_fill_1 FILLER_19_197 ();
 sg13g2_fill_2 FILLER_19_201 ();
 sg13g2_decap_4 FILLER_19_208 ();
 sg13g2_fill_2 FILLER_19_212 ();
 sg13g2_fill_1 FILLER_19_219 ();
 sg13g2_fill_2 FILLER_19_230 ();
 sg13g2_fill_1 FILLER_19_232 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_285 ();
 sg13g2_decap_4 FILLER_19_297 ();
 sg13g2_fill_2 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_352 ();
 sg13g2_fill_1 FILLER_19_372 ();
 sg13g2_decap_4 FILLER_19_378 ();
 sg13g2_fill_2 FILLER_19_382 ();
 sg13g2_fill_1 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_395 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_4 FILLER_19_409 ();
 sg13g2_fill_1 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_422 ();
 sg13g2_decap_4 FILLER_19_429 ();
 sg13g2_fill_2 FILLER_19_433 ();
 sg13g2_decap_4 FILLER_19_493 ();
 sg13g2_fill_1 FILLER_19_497 ();
 sg13g2_fill_2 FILLER_19_530 ();
 sg13g2_fill_1 FILLER_19_532 ();
 sg13g2_fill_2 FILLER_19_546 ();
 sg13g2_fill_1 FILLER_19_548 ();
 sg13g2_decap_8 FILLER_19_575 ();
 sg13g2_fill_1 FILLER_19_582 ();
 sg13g2_decap_4 FILLER_19_603 ();
 sg13g2_decap_4 FILLER_19_629 ();
 sg13g2_fill_1 FILLER_19_633 ();
 sg13g2_decap_8 FILLER_19_643 ();
 sg13g2_decap_4 FILLER_19_650 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_4 FILLER_19_693 ();
 sg13g2_fill_2 FILLER_19_697 ();
 sg13g2_fill_1 FILLER_19_727 ();
 sg13g2_decap_8 FILLER_19_746 ();
 sg13g2_decap_8 FILLER_19_753 ();
 sg13g2_decap_8 FILLER_19_760 ();
 sg13g2_fill_2 FILLER_19_767 ();
 sg13g2_fill_2 FILLER_19_795 ();
 sg13g2_fill_1 FILLER_19_797 ();
 sg13g2_fill_2 FILLER_19_812 ();
 sg13g2_decap_4 FILLER_19_823 ();
 sg13g2_decap_8 FILLER_19_837 ();
 sg13g2_fill_2 FILLER_19_844 ();
 sg13g2_fill_1 FILLER_19_846 ();
 sg13g2_fill_2 FILLER_19_862 ();
 sg13g2_fill_1 FILLER_19_864 ();
 sg13g2_fill_2 FILLER_19_885 ();
 sg13g2_fill_1 FILLER_19_907 ();
 sg13g2_decap_8 FILLER_19_920 ();
 sg13g2_decap_8 FILLER_19_927 ();
 sg13g2_decap_8 FILLER_19_959 ();
 sg13g2_decap_8 FILLER_19_966 ();
 sg13g2_decap_8 FILLER_19_973 ();
 sg13g2_decap_8 FILLER_19_980 ();
 sg13g2_decap_8 FILLER_19_987 ();
 sg13g2_decap_8 FILLER_19_994 ();
 sg13g2_decap_8 FILLER_19_1001 ();
 sg13g2_decap_8 FILLER_19_1008 ();
 sg13g2_decap_8 FILLER_19_1015 ();
 sg13g2_decap_8 FILLER_19_1022 ();
 sg13g2_fill_2 FILLER_20_4 ();
 sg13g2_decap_4 FILLER_20_10 ();
 sg13g2_fill_2 FILLER_20_14 ();
 sg13g2_decap_4 FILLER_20_38 ();
 sg13g2_fill_2 FILLER_20_42 ();
 sg13g2_fill_2 FILLER_20_70 ();
 sg13g2_fill_1 FILLER_20_72 ();
 sg13g2_decap_8 FILLER_20_90 ();
 sg13g2_decap_4 FILLER_20_97 ();
 sg13g2_fill_2 FILLER_20_101 ();
 sg13g2_fill_1 FILLER_20_116 ();
 sg13g2_decap_8 FILLER_20_131 ();
 sg13g2_decap_4 FILLER_20_161 ();
 sg13g2_fill_1 FILLER_20_165 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_4 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_221 ();
 sg13g2_decap_8 FILLER_20_228 ();
 sg13g2_decap_8 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_242 ();
 sg13g2_decap_8 FILLER_20_249 ();
 sg13g2_fill_2 FILLER_20_256 ();
 sg13g2_decap_4 FILLER_20_262 ();
 sg13g2_fill_2 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_fill_1 FILLER_20_280 ();
 sg13g2_fill_1 FILLER_20_295 ();
 sg13g2_fill_1 FILLER_20_345 ();
 sg13g2_fill_1 FILLER_20_359 ();
 sg13g2_fill_1 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_444 ();
 sg13g2_fill_1 FILLER_20_451 ();
 sg13g2_fill_2 FILLER_20_471 ();
 sg13g2_fill_2 FILLER_20_483 ();
 sg13g2_fill_1 FILLER_20_485 ();
 sg13g2_decap_8 FILLER_20_495 ();
 sg13g2_fill_1 FILLER_20_502 ();
 sg13g2_fill_2 FILLER_20_506 ();
 sg13g2_fill_2 FILLER_20_527 ();
 sg13g2_fill_1 FILLER_20_529 ();
 sg13g2_fill_1 FILLER_20_570 ();
 sg13g2_fill_2 FILLER_20_580 ();
 sg13g2_fill_1 FILLER_20_582 ();
 sg13g2_fill_1 FILLER_20_591 ();
 sg13g2_fill_2 FILLER_20_596 ();
 sg13g2_fill_1 FILLER_20_598 ();
 sg13g2_decap_8 FILLER_20_608 ();
 sg13g2_fill_2 FILLER_20_646 ();
 sg13g2_fill_1 FILLER_20_648 ();
 sg13g2_decap_4 FILLER_20_666 ();
 sg13g2_decap_8 FILLER_20_683 ();
 sg13g2_decap_8 FILLER_20_690 ();
 sg13g2_fill_1 FILLER_20_697 ();
 sg13g2_decap_4 FILLER_20_702 ();
 sg13g2_decap_8 FILLER_20_709 ();
 sg13g2_decap_8 FILLER_20_716 ();
 sg13g2_decap_4 FILLER_20_723 ();
 sg13g2_fill_1 FILLER_20_727 ();
 sg13g2_decap_4 FILLER_20_742 ();
 sg13g2_fill_1 FILLER_20_746 ();
 sg13g2_fill_1 FILLER_20_778 ();
 sg13g2_decap_4 FILLER_20_783 ();
 sg13g2_fill_2 FILLER_20_833 ();
 sg13g2_decap_8 FILLER_20_839 ();
 sg13g2_decap_8 FILLER_20_846 ();
 sg13g2_decap_8 FILLER_20_853 ();
 sg13g2_fill_1 FILLER_20_860 ();
 sg13g2_fill_2 FILLER_20_870 ();
 sg13g2_fill_1 FILLER_20_884 ();
 sg13g2_fill_1 FILLER_20_889 ();
 sg13g2_decap_8 FILLER_20_898 ();
 sg13g2_decap_8 FILLER_20_905 ();
 sg13g2_fill_2 FILLER_20_912 ();
 sg13g2_fill_1 FILLER_20_914 ();
 sg13g2_decap_4 FILLER_20_920 ();
 sg13g2_decap_8 FILLER_20_959 ();
 sg13g2_fill_1 FILLER_20_966 ();
 sg13g2_decap_8 FILLER_20_976 ();
 sg13g2_decap_8 FILLER_20_983 ();
 sg13g2_decap_8 FILLER_20_990 ();
 sg13g2_decap_8 FILLER_20_997 ();
 sg13g2_decap_8 FILLER_20_1004 ();
 sg13g2_decap_8 FILLER_20_1011 ();
 sg13g2_decap_8 FILLER_20_1018 ();
 sg13g2_decap_4 FILLER_20_1025 ();
 sg13g2_decap_8 FILLER_21_4 ();
 sg13g2_decap_4 FILLER_21_46 ();
 sg13g2_fill_1 FILLER_21_50 ();
 sg13g2_fill_2 FILLER_21_56 ();
 sg13g2_fill_1 FILLER_21_58 ();
 sg13g2_decap_8 FILLER_21_64 ();
 sg13g2_fill_2 FILLER_21_85 ();
 sg13g2_fill_1 FILLER_21_87 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_fill_1 FILLER_21_105 ();
 sg13g2_decap_4 FILLER_21_118 ();
 sg13g2_fill_1 FILLER_21_122 ();
 sg13g2_decap_8 FILLER_21_132 ();
 sg13g2_decap_8 FILLER_21_139 ();
 sg13g2_fill_2 FILLER_21_146 ();
 sg13g2_decap_4 FILLER_21_192 ();
 sg13g2_fill_2 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_202 ();
 sg13g2_fill_1 FILLER_21_222 ();
 sg13g2_fill_2 FILLER_21_233 ();
 sg13g2_fill_1 FILLER_21_235 ();
 sg13g2_fill_2 FILLER_21_276 ();
 sg13g2_decap_8 FILLER_21_309 ();
 sg13g2_fill_1 FILLER_21_316 ();
 sg13g2_decap_8 FILLER_21_352 ();
 sg13g2_fill_1 FILLER_21_359 ();
 sg13g2_fill_1 FILLER_21_392 ();
 sg13g2_fill_1 FILLER_21_397 ();
 sg13g2_decap_8 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_21_412 ();
 sg13g2_fill_2 FILLER_21_419 ();
 sg13g2_decap_4 FILLER_21_425 ();
 sg13g2_fill_2 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_21_444 ();
 sg13g2_decap_8 FILLER_21_451 ();
 sg13g2_decap_4 FILLER_21_458 ();
 sg13g2_fill_2 FILLER_21_462 ();
 sg13g2_decap_8 FILLER_21_491 ();
 sg13g2_decap_8 FILLER_21_526 ();
 sg13g2_fill_2 FILLER_21_533 ();
 sg13g2_fill_1 FILLER_21_535 ();
 sg13g2_fill_2 FILLER_21_549 ();
 sg13g2_fill_1 FILLER_21_551 ();
 sg13g2_decap_4 FILLER_21_562 ();
 sg13g2_decap_8 FILLER_21_575 ();
 sg13g2_decap_4 FILLER_21_582 ();
 sg13g2_decap_8 FILLER_21_614 ();
 sg13g2_decap_4 FILLER_21_621 ();
 sg13g2_fill_2 FILLER_21_625 ();
 sg13g2_decap_8 FILLER_21_633 ();
 sg13g2_decap_8 FILLER_21_640 ();
 sg13g2_fill_1 FILLER_21_647 ();
 sg13g2_fill_2 FILLER_21_661 ();
 sg13g2_decap_4 FILLER_21_667 ();
 sg13g2_fill_1 FILLER_21_671 ();
 sg13g2_decap_4 FILLER_21_685 ();
 sg13g2_fill_1 FILLER_21_689 ();
 sg13g2_fill_2 FILLER_21_726 ();
 sg13g2_fill_1 FILLER_21_728 ();
 sg13g2_decap_8 FILLER_21_777 ();
 sg13g2_decap_4 FILLER_21_784 ();
 sg13g2_fill_1 FILLER_21_788 ();
 sg13g2_fill_2 FILLER_21_793 ();
 sg13g2_fill_1 FILLER_21_799 ();
 sg13g2_decap_8 FILLER_21_816 ();
 sg13g2_fill_1 FILLER_21_823 ();
 sg13g2_decap_8 FILLER_21_843 ();
 sg13g2_fill_2 FILLER_21_850 ();
 sg13g2_fill_1 FILLER_21_852 ();
 sg13g2_fill_2 FILLER_21_866 ();
 sg13g2_fill_2 FILLER_21_886 ();
 sg13g2_fill_1 FILLER_21_888 ();
 sg13g2_fill_2 FILLER_21_894 ();
 sg13g2_decap_4 FILLER_21_909 ();
 sg13g2_fill_2 FILLER_21_913 ();
 sg13g2_decap_8 FILLER_21_920 ();
 sg13g2_decap_8 FILLER_21_927 ();
 sg13g2_fill_2 FILLER_21_934 ();
 sg13g2_fill_1 FILLER_21_954 ();
 sg13g2_decap_8 FILLER_21_983 ();
 sg13g2_decap_8 FILLER_21_990 ();
 sg13g2_decap_8 FILLER_21_997 ();
 sg13g2_decap_8 FILLER_21_1004 ();
 sg13g2_decap_8 FILLER_21_1011 ();
 sg13g2_decap_8 FILLER_21_1018 ();
 sg13g2_decap_4 FILLER_21_1025 ();
 sg13g2_fill_1 FILLER_22_43 ();
 sg13g2_fill_1 FILLER_22_49 ();
 sg13g2_fill_1 FILLER_22_53 ();
 sg13g2_decap_8 FILLER_22_58 ();
 sg13g2_fill_2 FILLER_22_65 ();
 sg13g2_fill_1 FILLER_22_89 ();
 sg13g2_fill_2 FILLER_22_106 ();
 sg13g2_decap_8 FILLER_22_136 ();
 sg13g2_decap_8 FILLER_22_143 ();
 sg13g2_decap_4 FILLER_22_150 ();
 sg13g2_fill_2 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_160 ();
 sg13g2_fill_1 FILLER_22_167 ();
 sg13g2_decap_4 FILLER_22_198 ();
 sg13g2_fill_1 FILLER_22_202 ();
 sg13g2_fill_2 FILLER_22_252 ();
 sg13g2_fill_1 FILLER_22_254 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_4 FILLER_22_280 ();
 sg13g2_decap_4 FILLER_22_288 ();
 sg13g2_fill_2 FILLER_22_292 ();
 sg13g2_decap_8 FILLER_22_303 ();
 sg13g2_fill_1 FILLER_22_310 ();
 sg13g2_fill_1 FILLER_22_377 ();
 sg13g2_decap_8 FILLER_22_404 ();
 sg13g2_decap_8 FILLER_22_411 ();
 sg13g2_decap_4 FILLER_22_418 ();
 sg13g2_fill_2 FILLER_22_422 ();
 sg13g2_fill_2 FILLER_22_427 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_4 FILLER_22_434 ();
 sg13g2_fill_1 FILLER_22_438 ();
 sg13g2_decap_8 FILLER_22_452 ();
 sg13g2_decap_4 FILLER_22_459 ();
 sg13g2_decap_4 FILLER_22_485 ();
 sg13g2_fill_1 FILLER_22_489 ();
 sg13g2_decap_8 FILLER_22_507 ();
 sg13g2_decap_8 FILLER_22_514 ();
 sg13g2_decap_8 FILLER_22_521 ();
 sg13g2_decap_4 FILLER_22_528 ();
 sg13g2_fill_1 FILLER_22_545 ();
 sg13g2_fill_2 FILLER_22_577 ();
 sg13g2_decap_8 FILLER_22_622 ();
 sg13g2_decap_8 FILLER_22_629 ();
 sg13g2_fill_2 FILLER_22_636 ();
 sg13g2_fill_1 FILLER_22_638 ();
 sg13g2_decap_8 FILLER_22_643 ();
 sg13g2_decap_8 FILLER_22_650 ();
 sg13g2_fill_1 FILLER_22_657 ();
 sg13g2_fill_1 FILLER_22_714 ();
 sg13g2_decap_8 FILLER_22_739 ();
 sg13g2_fill_1 FILLER_22_746 ();
 sg13g2_fill_2 FILLER_22_757 ();
 sg13g2_decap_4 FILLER_22_764 ();
 sg13g2_fill_1 FILLER_22_768 ();
 sg13g2_decap_4 FILLER_22_778 ();
 sg13g2_fill_2 FILLER_22_782 ();
 sg13g2_decap_8 FILLER_22_815 ();
 sg13g2_fill_2 FILLER_22_822 ();
 sg13g2_fill_1 FILLER_22_824 ();
 sg13g2_fill_2 FILLER_22_880 ();
 sg13g2_fill_1 FILLER_22_882 ();
 sg13g2_fill_2 FILLER_22_892 ();
 sg13g2_decap_8 FILLER_22_907 ();
 sg13g2_fill_2 FILLER_22_914 ();
 sg13g2_fill_2 FILLER_22_920 ();
 sg13g2_decap_8 FILLER_22_935 ();
 sg13g2_fill_2 FILLER_22_942 ();
 sg13g2_fill_1 FILLER_22_944 ();
 sg13g2_decap_8 FILLER_22_950 ();
 sg13g2_fill_2 FILLER_22_957 ();
 sg13g2_fill_1 FILLER_22_959 ();
 sg13g2_decap_8 FILLER_22_964 ();
 sg13g2_decap_8 FILLER_22_971 ();
 sg13g2_decap_8 FILLER_22_978 ();
 sg13g2_decap_8 FILLER_22_985 ();
 sg13g2_decap_8 FILLER_22_992 ();
 sg13g2_decap_8 FILLER_22_999 ();
 sg13g2_decap_8 FILLER_22_1006 ();
 sg13g2_decap_8 FILLER_22_1013 ();
 sg13g2_decap_8 FILLER_22_1020 ();
 sg13g2_fill_2 FILLER_22_1027 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_41 ();
 sg13g2_fill_1 FILLER_23_52 ();
 sg13g2_decap_4 FILLER_23_63 ();
 sg13g2_fill_2 FILLER_23_67 ();
 sg13g2_decap_8 FILLER_23_101 ();
 sg13g2_decap_8 FILLER_23_108 ();
 sg13g2_decap_4 FILLER_23_128 ();
 sg13g2_decap_8 FILLER_23_159 ();
 sg13g2_decap_4 FILLER_23_179 ();
 sg13g2_fill_2 FILLER_23_193 ();
 sg13g2_fill_1 FILLER_23_195 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_fill_2 FILLER_23_224 ();
 sg13g2_fill_1 FILLER_23_239 ();
 sg13g2_decap_4 FILLER_23_262 ();
 sg13g2_fill_2 FILLER_23_276 ();
 sg13g2_fill_1 FILLER_23_278 ();
 sg13g2_fill_2 FILLER_23_335 ();
 sg13g2_decap_8 FILLER_23_341 ();
 sg13g2_decap_8 FILLER_23_365 ();
 sg13g2_decap_4 FILLER_23_372 ();
 sg13g2_fill_1 FILLER_23_466 ();
 sg13g2_decap_8 FILLER_23_480 ();
 sg13g2_decap_8 FILLER_23_487 ();
 sg13g2_decap_8 FILLER_23_494 ();
 sg13g2_decap_8 FILLER_23_501 ();
 sg13g2_fill_1 FILLER_23_508 ();
 sg13g2_fill_2 FILLER_23_537 ();
 sg13g2_fill_1 FILLER_23_539 ();
 sg13g2_fill_2 FILLER_23_553 ();
 sg13g2_fill_2 FILLER_23_559 ();
 sg13g2_fill_2 FILLER_23_565 ();
 sg13g2_fill_1 FILLER_23_567 ();
 sg13g2_decap_4 FILLER_23_577 ();
 sg13g2_fill_1 FILLER_23_581 ();
 sg13g2_decap_4 FILLER_23_669 ();
 sg13g2_fill_1 FILLER_23_702 ();
 sg13g2_fill_1 FILLER_23_737 ();
 sg13g2_fill_2 FILLER_23_773 ();
 sg13g2_fill_2 FILLER_23_790 ();
 sg13g2_fill_2 FILLER_23_814 ();
 sg13g2_decap_8 FILLER_23_835 ();
 sg13g2_decap_8 FILLER_23_842 ();
 sg13g2_decap_8 FILLER_23_849 ();
 sg13g2_fill_1 FILLER_23_856 ();
 sg13g2_decap_4 FILLER_23_861 ();
 sg13g2_fill_2 FILLER_23_865 ();
 sg13g2_decap_8 FILLER_23_871 ();
 sg13g2_fill_2 FILLER_23_878 ();
 sg13g2_fill_2 FILLER_23_907 ();
 sg13g2_fill_1 FILLER_23_909 ();
 sg13g2_decap_8 FILLER_23_950 ();
 sg13g2_decap_8 FILLER_23_957 ();
 sg13g2_decap_8 FILLER_23_964 ();
 sg13g2_decap_8 FILLER_23_971 ();
 sg13g2_decap_8 FILLER_23_978 ();
 sg13g2_decap_8 FILLER_23_985 ();
 sg13g2_decap_8 FILLER_23_992 ();
 sg13g2_decap_8 FILLER_23_999 ();
 sg13g2_decap_8 FILLER_23_1006 ();
 sg13g2_decap_8 FILLER_23_1013 ();
 sg13g2_decap_8 FILLER_23_1020 ();
 sg13g2_fill_2 FILLER_23_1027 ();
 sg13g2_fill_2 FILLER_24_4 ();
 sg13g2_decap_8 FILLER_24_10 ();
 sg13g2_decap_4 FILLER_24_17 ();
 sg13g2_fill_2 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_66 ();
 sg13g2_fill_2 FILLER_24_73 ();
 sg13g2_decap_4 FILLER_24_83 ();
 sg13g2_fill_1 FILLER_24_87 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_4 FILLER_24_112 ();
 sg13g2_decap_4 FILLER_24_143 ();
 sg13g2_fill_2 FILLER_24_160 ();
 sg13g2_fill_1 FILLER_24_162 ();
 sg13g2_decap_4 FILLER_24_172 ();
 sg13g2_fill_2 FILLER_24_176 ();
 sg13g2_fill_2 FILLER_24_191 ();
 sg13g2_fill_1 FILLER_24_193 ();
 sg13g2_fill_1 FILLER_24_221 ();
 sg13g2_decap_8 FILLER_24_258 ();
 sg13g2_fill_1 FILLER_24_278 ();
 sg13g2_decap_8 FILLER_24_288 ();
 sg13g2_decap_4 FILLER_24_295 ();
 sg13g2_decap_8 FILLER_24_321 ();
 sg13g2_decap_4 FILLER_24_328 ();
 sg13g2_fill_1 FILLER_24_335 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_fill_2 FILLER_24_371 ();
 sg13g2_fill_1 FILLER_24_373 ();
 sg13g2_fill_2 FILLER_24_397 ();
 sg13g2_fill_1 FILLER_24_399 ();
 sg13g2_decap_8 FILLER_24_434 ();
 sg13g2_fill_2 FILLER_24_450 ();
 sg13g2_fill_1 FILLER_24_452 ();
 sg13g2_decap_8 FILLER_24_468 ();
 sg13g2_decap_4 FILLER_24_475 ();
 sg13g2_fill_2 FILLER_24_479 ();
 sg13g2_fill_1 FILLER_24_496 ();
 sg13g2_fill_1 FILLER_24_509 ();
 sg13g2_decap_8 FILLER_24_527 ();
 sg13g2_decap_8 FILLER_24_534 ();
 sg13g2_decap_8 FILLER_24_541 ();
 sg13g2_decap_8 FILLER_24_591 ();
 sg13g2_decap_8 FILLER_24_598 ();
 sg13g2_decap_4 FILLER_24_605 ();
 sg13g2_decap_8 FILLER_24_617 ();
 sg13g2_fill_2 FILLER_24_624 ();
 sg13g2_decap_4 FILLER_24_643 ();
 sg13g2_fill_2 FILLER_24_647 ();
 sg13g2_decap_8 FILLER_24_676 ();
 sg13g2_fill_2 FILLER_24_711 ();
 sg13g2_fill_1 FILLER_24_713 ();
 sg13g2_fill_2 FILLER_24_734 ();
 sg13g2_fill_1 FILLER_24_736 ();
 sg13g2_fill_2 FILLER_24_742 ();
 sg13g2_fill_2 FILLER_24_752 ();
 sg13g2_fill_2 FILLER_24_759 ();
 sg13g2_decap_8 FILLER_24_766 ();
 sg13g2_decap_4 FILLER_24_773 ();
 sg13g2_fill_2 FILLER_24_777 ();
 sg13g2_decap_8 FILLER_24_812 ();
 sg13g2_fill_2 FILLER_24_819 ();
 sg13g2_fill_1 FILLER_24_821 ();
 sg13g2_decap_8 FILLER_24_835 ();
 sg13g2_fill_1 FILLER_24_842 ();
 sg13g2_fill_1 FILLER_24_870 ();
 sg13g2_decap_8 FILLER_24_875 ();
 sg13g2_decap_4 FILLER_24_887 ();
 sg13g2_fill_2 FILLER_24_891 ();
 sg13g2_fill_1 FILLER_24_903 ();
 sg13g2_fill_1 FILLER_24_917 ();
 sg13g2_fill_2 FILLER_24_923 ();
 sg13g2_decap_8 FILLER_24_965 ();
 sg13g2_decap_8 FILLER_24_972 ();
 sg13g2_decap_8 FILLER_24_979 ();
 sg13g2_decap_8 FILLER_24_986 ();
 sg13g2_decap_8 FILLER_24_993 ();
 sg13g2_decap_8 FILLER_24_1000 ();
 sg13g2_decap_8 FILLER_24_1007 ();
 sg13g2_decap_8 FILLER_24_1014 ();
 sg13g2_decap_8 FILLER_24_1021 ();
 sg13g2_fill_1 FILLER_24_1028 ();
 sg13g2_decap_8 FILLER_25_4 ();
 sg13g2_decap_8 FILLER_25_11 ();
 sg13g2_decap_8 FILLER_25_18 ();
 sg13g2_decap_8 FILLER_25_25 ();
 sg13g2_fill_2 FILLER_25_32 ();
 sg13g2_fill_1 FILLER_25_34 ();
 sg13g2_fill_1 FILLER_25_39 ();
 sg13g2_decap_4 FILLER_25_45 ();
 sg13g2_fill_1 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_132 ();
 sg13g2_decap_8 FILLER_25_139 ();
 sg13g2_decap_4 FILLER_25_146 ();
 sg13g2_fill_1 FILLER_25_150 ();
 sg13g2_fill_2 FILLER_25_182 ();
 sg13g2_fill_1 FILLER_25_184 ();
 sg13g2_decap_8 FILLER_25_213 ();
 sg13g2_fill_2 FILLER_25_234 ();
 sg13g2_fill_1 FILLER_25_240 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_fill_2 FILLER_25_252 ();
 sg13g2_fill_1 FILLER_25_254 ();
 sg13g2_decap_8 FILLER_25_290 ();
 sg13g2_decap_4 FILLER_25_297 ();
 sg13g2_fill_2 FILLER_25_316 ();
 sg13g2_decap_8 FILLER_25_332 ();
 sg13g2_fill_2 FILLER_25_339 ();
 sg13g2_fill_1 FILLER_25_345 ();
 sg13g2_decap_8 FILLER_25_355 ();
 sg13g2_decap_4 FILLER_25_362 ();
 sg13g2_fill_1 FILLER_25_366 ();
 sg13g2_decap_4 FILLER_25_380 ();
 sg13g2_fill_2 FILLER_25_384 ();
 sg13g2_fill_1 FILLER_25_406 ();
 sg13g2_fill_2 FILLER_25_431 ();
 sg13g2_fill_1 FILLER_25_433 ();
 sg13g2_decap_4 FILLER_25_444 ();
 sg13g2_fill_1 FILLER_25_448 ();
 sg13g2_fill_2 FILLER_25_464 ();
 sg13g2_fill_1 FILLER_25_466 ();
 sg13g2_decap_4 FILLER_25_538 ();
 sg13g2_decap_8 FILLER_25_562 ();
 sg13g2_fill_2 FILLER_25_569 ();
 sg13g2_fill_1 FILLER_25_571 ();
 sg13g2_decap_8 FILLER_25_587 ();
 sg13g2_fill_1 FILLER_25_594 ();
 sg13g2_decap_4 FILLER_25_623 ();
 sg13g2_fill_2 FILLER_25_627 ();
 sg13g2_fill_1 FILLER_25_648 ();
 sg13g2_decap_4 FILLER_25_679 ();
 sg13g2_decap_4 FILLER_25_695 ();
 sg13g2_fill_2 FILLER_25_699 ();
 sg13g2_fill_2 FILLER_25_710 ();
 sg13g2_fill_1 FILLER_25_712 ();
 sg13g2_decap_8 FILLER_25_733 ();
 sg13g2_decap_8 FILLER_25_740 ();
 sg13g2_decap_8 FILLER_25_747 ();
 sg13g2_fill_1 FILLER_25_763 ();
 sg13g2_decap_8 FILLER_25_768 ();
 sg13g2_fill_2 FILLER_25_775 ();
 sg13g2_decap_4 FILLER_25_808 ();
 sg13g2_fill_2 FILLER_25_843 ();
 sg13g2_fill_1 FILLER_25_845 ();
 sg13g2_decap_4 FILLER_25_860 ();
 sg13g2_fill_2 FILLER_25_864 ();
 sg13g2_decap_8 FILLER_25_894 ();
 sg13g2_fill_2 FILLER_25_901 ();
 sg13g2_fill_2 FILLER_25_914 ();
 sg13g2_decap_4 FILLER_25_926 ();
 sg13g2_fill_2 FILLER_25_930 ();
 sg13g2_decap_8 FILLER_25_985 ();
 sg13g2_decap_8 FILLER_25_992 ();
 sg13g2_decap_8 FILLER_25_999 ();
 sg13g2_decap_8 FILLER_25_1006 ();
 sg13g2_decap_8 FILLER_25_1013 ();
 sg13g2_decap_8 FILLER_25_1020 ();
 sg13g2_fill_2 FILLER_25_1027 ();
 sg13g2_decap_8 FILLER_26_4 ();
 sg13g2_decap_8 FILLER_26_15 ();
 sg13g2_decap_8 FILLER_26_22 ();
 sg13g2_decap_8 FILLER_26_29 ();
 sg13g2_fill_1 FILLER_26_36 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_4 FILLER_26_56 ();
 sg13g2_fill_2 FILLER_26_60 ();
 sg13g2_decap_8 FILLER_26_79 ();
 sg13g2_decap_8 FILLER_26_86 ();
 sg13g2_decap_8 FILLER_26_93 ();
 sg13g2_decap_4 FILLER_26_100 ();
 sg13g2_decap_8 FILLER_26_178 ();
 sg13g2_decap_4 FILLER_26_185 ();
 sg13g2_fill_1 FILLER_26_189 ();
 sg13g2_fill_2 FILLER_26_202 ();
 sg13g2_fill_1 FILLER_26_204 ();
 sg13g2_decap_4 FILLER_26_214 ();
 sg13g2_fill_2 FILLER_26_218 ();
 sg13g2_decap_8 FILLER_26_240 ();
 sg13g2_decap_8 FILLER_26_247 ();
 sg13g2_fill_1 FILLER_26_254 ();
 sg13g2_decap_8 FILLER_26_270 ();
 sg13g2_fill_1 FILLER_26_277 ();
 sg13g2_decap_4 FILLER_26_287 ();
 sg13g2_fill_2 FILLER_26_311 ();
 sg13g2_fill_2 FILLER_26_318 ();
 sg13g2_decap_8 FILLER_26_337 ();
 sg13g2_fill_1 FILLER_26_347 ();
 sg13g2_fill_2 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_406 ();
 sg13g2_fill_2 FILLER_26_413 ();
 sg13g2_fill_1 FILLER_26_415 ();
 sg13g2_decap_8 FILLER_26_434 ();
 sg13g2_decap_8 FILLER_26_441 ();
 sg13g2_decap_8 FILLER_26_448 ();
 sg13g2_fill_1 FILLER_26_470 ();
 sg13g2_fill_1 FILLER_26_479 ();
 sg13g2_decap_8 FILLER_26_495 ();
 sg13g2_fill_1 FILLER_26_502 ();
 sg13g2_decap_8 FILLER_26_508 ();
 sg13g2_decap_4 FILLER_26_515 ();
 sg13g2_fill_2 FILLER_26_519 ();
 sg13g2_decap_4 FILLER_26_530 ();
 sg13g2_fill_2 FILLER_26_534 ();
 sg13g2_decap_8 FILLER_26_561 ();
 sg13g2_fill_2 FILLER_26_568 ();
 sg13g2_decap_4 FILLER_26_590 ();
 sg13g2_fill_1 FILLER_26_594 ();
 sg13g2_decap_8 FILLER_26_640 ();
 sg13g2_decap_8 FILLER_26_647 ();
 sg13g2_fill_2 FILLER_26_654 ();
 sg13g2_fill_1 FILLER_26_656 ();
 sg13g2_decap_8 FILLER_26_681 ();
 sg13g2_fill_2 FILLER_26_688 ();
 sg13g2_fill_1 FILLER_26_694 ();
 sg13g2_decap_8 FILLER_26_700 ();
 sg13g2_fill_1 FILLER_26_707 ();
 sg13g2_decap_4 FILLER_26_713 ();
 sg13g2_decap_8 FILLER_26_727 ();
 sg13g2_fill_2 FILLER_26_734 ();
 sg13g2_decap_4 FILLER_26_740 ();
 sg13g2_decap_8 FILLER_26_749 ();
 sg13g2_fill_1 FILLER_26_756 ();
 sg13g2_decap_4 FILLER_26_778 ();
 sg13g2_decap_8 FILLER_26_797 ();
 sg13g2_decap_4 FILLER_26_804 ();
 sg13g2_fill_1 FILLER_26_827 ();
 sg13g2_decap_8 FILLER_26_852 ();
 sg13g2_decap_4 FILLER_26_859 ();
 sg13g2_fill_2 FILLER_26_863 ();
 sg13g2_decap_8 FILLER_26_878 ();
 sg13g2_decap_8 FILLER_26_885 ();
 sg13g2_decap_8 FILLER_26_892 ();
 sg13g2_fill_2 FILLER_26_899 ();
 sg13g2_decap_4 FILLER_26_926 ();
 sg13g2_fill_1 FILLER_26_930 ();
 sg13g2_fill_2 FILLER_26_948 ();
 sg13g2_fill_1 FILLER_26_950 ();
 sg13g2_fill_2 FILLER_26_961 ();
 sg13g2_decap_4 FILLER_26_967 ();
 sg13g2_decap_8 FILLER_26_980 ();
 sg13g2_decap_8 FILLER_26_987 ();
 sg13g2_decap_8 FILLER_26_994 ();
 sg13g2_decap_8 FILLER_26_1001 ();
 sg13g2_decap_8 FILLER_26_1008 ();
 sg13g2_decap_8 FILLER_26_1015 ();
 sg13g2_decap_8 FILLER_26_1022 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_4 ();
 sg13g2_fill_1 FILLER_27_41 ();
 sg13g2_decap_8 FILLER_27_52 ();
 sg13g2_fill_2 FILLER_27_59 ();
 sg13g2_fill_1 FILLER_27_61 ();
 sg13g2_fill_2 FILLER_27_82 ();
 sg13g2_fill_1 FILLER_27_84 ();
 sg13g2_fill_2 FILLER_27_94 ();
 sg13g2_fill_1 FILLER_27_96 ();
 sg13g2_fill_2 FILLER_27_112 ();
 sg13g2_fill_2 FILLER_27_119 ();
 sg13g2_decap_4 FILLER_27_183 ();
 sg13g2_fill_1 FILLER_27_187 ();
 sg13g2_fill_2 FILLER_27_195 ();
 sg13g2_decap_8 FILLER_27_201 ();
 sg13g2_fill_1 FILLER_27_221 ();
 sg13g2_fill_2 FILLER_27_237 ();
 sg13g2_fill_2 FILLER_27_244 ();
 sg13g2_decap_8 FILLER_27_275 ();
 sg13g2_decap_8 FILLER_27_282 ();
 sg13g2_fill_2 FILLER_27_289 ();
 sg13g2_fill_1 FILLER_27_291 ();
 sg13g2_fill_2 FILLER_27_302 ();
 sg13g2_fill_2 FILLER_27_314 ();
 sg13g2_fill_1 FILLER_27_316 ();
 sg13g2_fill_1 FILLER_27_322 ();
 sg13g2_decap_4 FILLER_27_333 ();
 sg13g2_decap_4 FILLER_27_342 ();
 sg13g2_fill_2 FILLER_27_346 ();
 sg13g2_fill_2 FILLER_27_370 ();
 sg13g2_fill_1 FILLER_27_372 ();
 sg13g2_fill_1 FILLER_27_377 ();
 sg13g2_decap_8 FILLER_27_382 ();
 sg13g2_fill_2 FILLER_27_389 ();
 sg13g2_fill_1 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_409 ();
 sg13g2_fill_2 FILLER_27_416 ();
 sg13g2_decap_8 FILLER_27_433 ();
 sg13g2_decap_8 FILLER_27_440 ();
 sg13g2_decap_8 FILLER_27_447 ();
 sg13g2_decap_8 FILLER_27_454 ();
 sg13g2_decap_4 FILLER_27_461 ();
 sg13g2_decap_4 FILLER_27_484 ();
 sg13g2_decap_4 FILLER_27_493 ();
 sg13g2_fill_1 FILLER_27_497 ();
 sg13g2_decap_4 FILLER_27_501 ();
 sg13g2_fill_2 FILLER_27_505 ();
 sg13g2_fill_1 FILLER_27_511 ();
 sg13g2_decap_8 FILLER_27_529 ();
 sg13g2_decap_8 FILLER_27_536 ();
 sg13g2_decap_4 FILLER_27_543 ();
 sg13g2_fill_1 FILLER_27_547 ();
 sg13g2_decap_4 FILLER_27_557 ();
 sg13g2_fill_2 FILLER_27_561 ();
 sg13g2_fill_2 FILLER_27_568 ();
 sg13g2_fill_1 FILLER_27_570 ();
 sg13g2_decap_8 FILLER_27_585 ();
 sg13g2_decap_8 FILLER_27_592 ();
 sg13g2_decap_8 FILLER_27_599 ();
 sg13g2_fill_1 FILLER_27_606 ();
 sg13g2_fill_1 FILLER_27_625 ();
 sg13g2_decap_8 FILLER_27_643 ();
 sg13g2_decap_8 FILLER_27_650 ();
 sg13g2_fill_1 FILLER_27_670 ();
 sg13g2_fill_2 FILLER_27_676 ();
 sg13g2_decap_8 FILLER_27_703 ();
 sg13g2_decap_8 FILLER_27_710 ();
 sg13g2_decap_8 FILLER_27_717 ();
 sg13g2_fill_2 FILLER_27_724 ();
 sg13g2_fill_1 FILLER_27_726 ();
 sg13g2_fill_1 FILLER_27_737 ();
 sg13g2_fill_2 FILLER_27_742 ();
 sg13g2_fill_1 FILLER_27_744 ();
 sg13g2_decap_8 FILLER_27_753 ();
 sg13g2_fill_2 FILLER_27_760 ();
 sg13g2_decap_8 FILLER_27_767 ();
 sg13g2_decap_4 FILLER_27_774 ();
 sg13g2_fill_1 FILLER_27_778 ();
 sg13g2_decap_4 FILLER_27_784 ();
 sg13g2_fill_1 FILLER_27_800 ();
 sg13g2_decap_8 FILLER_27_806 ();
 sg13g2_decap_4 FILLER_27_813 ();
 sg13g2_fill_1 FILLER_27_817 ();
 sg13g2_decap_4 FILLER_27_835 ();
 sg13g2_decap_8 FILLER_27_851 ();
 sg13g2_decap_8 FILLER_27_858 ();
 sg13g2_decap_4 FILLER_27_865 ();
 sg13g2_fill_2 FILLER_27_869 ();
 sg13g2_decap_8 FILLER_27_885 ();
 sg13g2_fill_2 FILLER_27_892 ();
 sg13g2_fill_1 FILLER_27_894 ();
 sg13g2_decap_8 FILLER_27_918 ();
 sg13g2_fill_1 FILLER_27_925 ();
 sg13g2_fill_1 FILLER_27_956 ();
 sg13g2_decap_8 FILLER_27_988 ();
 sg13g2_decap_8 FILLER_27_995 ();
 sg13g2_decap_8 FILLER_27_1002 ();
 sg13g2_decap_8 FILLER_27_1009 ();
 sg13g2_decap_8 FILLER_27_1016 ();
 sg13g2_decap_4 FILLER_27_1023 ();
 sg13g2_fill_2 FILLER_27_1027 ();
 sg13g2_decap_4 FILLER_28_4 ();
 sg13g2_decap_4 FILLER_28_15 ();
 sg13g2_fill_2 FILLER_28_19 ();
 sg13g2_decap_4 FILLER_28_45 ();
 sg13g2_fill_1 FILLER_28_85 ();
 sg13g2_fill_2 FILLER_28_91 ();
 sg13g2_fill_1 FILLER_28_93 ();
 sg13g2_fill_1 FILLER_28_109 ();
 sg13g2_fill_1 FILLER_28_126 ();
 sg13g2_fill_2 FILLER_28_131 ();
 sg13g2_fill_2 FILLER_28_148 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_265 ();
 sg13g2_decap_8 FILLER_28_272 ();
 sg13g2_fill_2 FILLER_28_279 ();
 sg13g2_fill_1 FILLER_28_281 ();
 sg13g2_fill_2 FILLER_28_295 ();
 sg13g2_decap_4 FILLER_28_317 ();
 sg13g2_fill_2 FILLER_28_321 ();
 sg13g2_fill_1 FILLER_28_328 ();
 sg13g2_decap_8 FILLER_28_339 ();
 sg13g2_decap_8 FILLER_28_346 ();
 sg13g2_fill_2 FILLER_28_357 ();
 sg13g2_fill_1 FILLER_28_372 ();
 sg13g2_fill_2 FILLER_28_439 ();
 sg13g2_decap_8 FILLER_28_446 ();
 sg13g2_fill_1 FILLER_28_453 ();
 sg13g2_fill_1 FILLER_28_459 ();
 sg13g2_fill_2 FILLER_28_477 ();
 sg13g2_fill_1 FILLER_28_479 ();
 sg13g2_fill_2 FILLER_28_486 ();
 sg13g2_decap_8 FILLER_28_558 ();
 sg13g2_fill_2 FILLER_28_565 ();
 sg13g2_decap_8 FILLER_28_590 ();
 sg13g2_decap_8 FILLER_28_597 ();
 sg13g2_fill_2 FILLER_28_604 ();
 sg13g2_fill_1 FILLER_28_611 ();
 sg13g2_fill_2 FILLER_28_617 ();
 sg13g2_fill_1 FILLER_28_619 ();
 sg13g2_fill_2 FILLER_28_625 ();
 sg13g2_decap_8 FILLER_28_638 ();
 sg13g2_decap_8 FILLER_28_645 ();
 sg13g2_fill_2 FILLER_28_652 ();
 sg13g2_decap_8 FILLER_28_667 ();
 sg13g2_fill_2 FILLER_28_674 ();
 sg13g2_fill_1 FILLER_28_676 ();
 sg13g2_decap_8 FILLER_28_705 ();
 sg13g2_fill_1 FILLER_28_712 ();
 sg13g2_fill_2 FILLER_28_718 ();
 sg13g2_fill_1 FILLER_28_720 ();
 sg13g2_fill_2 FILLER_28_756 ();
 sg13g2_decap_4 FILLER_28_782 ();
 sg13g2_decap_8 FILLER_28_795 ();
 sg13g2_fill_1 FILLER_28_802 ();
 sg13g2_fill_1 FILLER_28_806 ();
 sg13g2_fill_1 FILLER_28_835 ();
 sg13g2_fill_1 FILLER_28_844 ();
 sg13g2_fill_1 FILLER_28_861 ();
 sg13g2_decap_4 FILLER_28_889 ();
 sg13g2_fill_1 FILLER_28_893 ();
 sg13g2_decap_8 FILLER_28_909 ();
 sg13g2_decap_8 FILLER_28_916 ();
 sg13g2_decap_4 FILLER_28_923 ();
 sg13g2_fill_1 FILLER_28_927 ();
 sg13g2_fill_1 FILLER_28_948 ();
 sg13g2_decap_8 FILLER_28_954 ();
 sg13g2_decap_4 FILLER_28_961 ();
 sg13g2_fill_1 FILLER_28_969 ();
 sg13g2_decap_8 FILLER_28_979 ();
 sg13g2_decap_8 FILLER_28_986 ();
 sg13g2_decap_8 FILLER_28_993 ();
 sg13g2_decap_8 FILLER_28_1000 ();
 sg13g2_decap_8 FILLER_28_1007 ();
 sg13g2_decap_8 FILLER_28_1014 ();
 sg13g2_decap_8 FILLER_28_1021 ();
 sg13g2_fill_1 FILLER_28_1028 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_1 FILLER_29_31 ();
 sg13g2_fill_2 FILLER_29_41 ();
 sg13g2_fill_2 FILLER_29_56 ();
 sg13g2_fill_1 FILLER_29_58 ();
 sg13g2_fill_1 FILLER_29_88 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_fill_1 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_151 ();
 sg13g2_fill_1 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_181 ();
 sg13g2_decap_8 FILLER_29_188 ();
 sg13g2_decap_8 FILLER_29_195 ();
 sg13g2_decap_8 FILLER_29_211 ();
 sg13g2_fill_2 FILLER_29_218 ();
 sg13g2_decap_8 FILLER_29_238 ();
 sg13g2_fill_1 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_decap_4 FILLER_29_266 ();
 sg13g2_fill_2 FILLER_29_270 ();
 sg13g2_decap_8 FILLER_29_285 ();
 sg13g2_fill_2 FILLER_29_292 ();
 sg13g2_fill_2 FILLER_29_304 ();
 sg13g2_fill_1 FILLER_29_306 ();
 sg13g2_decap_4 FILLER_29_314 ();
 sg13g2_fill_1 FILLER_29_334 ();
 sg13g2_fill_2 FILLER_29_340 ();
 sg13g2_fill_2 FILLER_29_345 ();
 sg13g2_fill_2 FILLER_29_375 ();
 sg13g2_fill_1 FILLER_29_377 ();
 sg13g2_decap_8 FILLER_29_381 ();
 sg13g2_decap_8 FILLER_29_388 ();
 sg13g2_decap_8 FILLER_29_395 ();
 sg13g2_fill_2 FILLER_29_402 ();
 sg13g2_fill_2 FILLER_29_418 ();
 sg13g2_fill_1 FILLER_29_420 ();
 sg13g2_decap_8 FILLER_29_435 ();
 sg13g2_decap_8 FILLER_29_442 ();
 sg13g2_fill_2 FILLER_29_449 ();
 sg13g2_fill_1 FILLER_29_451 ();
 sg13g2_decap_8 FILLER_29_492 ();
 sg13g2_decap_8 FILLER_29_499 ();
 sg13g2_decap_4 FILLER_29_506 ();
 sg13g2_fill_2 FILLER_29_510 ();
 sg13g2_fill_2 FILLER_29_521 ();
 sg13g2_fill_1 FILLER_29_523 ();
 sg13g2_decap_8 FILLER_29_533 ();
 sg13g2_fill_1 FILLER_29_540 ();
 sg13g2_decap_4 FILLER_29_561 ();
 sg13g2_fill_2 FILLER_29_565 ();
 sg13g2_fill_2 FILLER_29_577 ();
 sg13g2_decap_8 FILLER_29_584 ();
 sg13g2_fill_1 FILLER_29_591 ();
 sg13g2_decap_8 FILLER_29_596 ();
 sg13g2_decap_8 FILLER_29_638 ();
 sg13g2_fill_1 FILLER_29_650 ();
 sg13g2_fill_1 FILLER_29_656 ();
 sg13g2_fill_1 FILLER_29_661 ();
 sg13g2_fill_2 FILLER_29_681 ();
 sg13g2_fill_1 FILLER_29_683 ();
 sg13g2_decap_8 FILLER_29_699 ();
 sg13g2_fill_2 FILLER_29_706 ();
 sg13g2_decap_8 FILLER_29_712 ();
 sg13g2_decap_8 FILLER_29_719 ();
 sg13g2_fill_1 FILLER_29_731 ();
 sg13g2_fill_1 FILLER_29_763 ();
 sg13g2_decap_8 FILLER_29_769 ();
 sg13g2_fill_2 FILLER_29_776 ();
 sg13g2_decap_4 FILLER_29_808 ();
 sg13g2_fill_1 FILLER_29_816 ();
 sg13g2_decap_8 FILLER_29_829 ();
 sg13g2_decap_8 FILLER_29_836 ();
 sg13g2_fill_2 FILLER_29_843 ();
 sg13g2_decap_8 FILLER_29_855 ();
 sg13g2_decap_8 FILLER_29_862 ();
 sg13g2_fill_2 FILLER_29_869 ();
 sg13g2_decap_8 FILLER_29_881 ();
 sg13g2_fill_1 FILLER_29_888 ();
 sg13g2_fill_2 FILLER_29_903 ();
 sg13g2_fill_1 FILLER_29_905 ();
 sg13g2_decap_4 FILLER_29_919 ();
 sg13g2_fill_2 FILLER_29_923 ();
 sg13g2_fill_1 FILLER_29_930 ();
 sg13g2_fill_2 FILLER_29_936 ();
 sg13g2_fill_1 FILLER_29_957 ();
 sg13g2_fill_2 FILLER_29_962 ();
 sg13g2_fill_1 FILLER_29_964 ();
 sg13g2_decap_8 FILLER_29_974 ();
 sg13g2_decap_8 FILLER_29_981 ();
 sg13g2_decap_8 FILLER_29_988 ();
 sg13g2_decap_8 FILLER_29_995 ();
 sg13g2_decap_8 FILLER_29_1002 ();
 sg13g2_decap_8 FILLER_29_1009 ();
 sg13g2_decap_8 FILLER_29_1016 ();
 sg13g2_decap_4 FILLER_29_1023 ();
 sg13g2_fill_2 FILLER_29_1027 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_9 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_4 FILLER_30_28 ();
 sg13g2_fill_1 FILLER_30_32 ();
 sg13g2_fill_2 FILLER_30_51 ();
 sg13g2_fill_1 FILLER_30_53 ();
 sg13g2_fill_1 FILLER_30_63 ();
 sg13g2_fill_1 FILLER_30_74 ();
 sg13g2_decap_8 FILLER_30_93 ();
 sg13g2_fill_2 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_118 ();
 sg13g2_decap_8 FILLER_30_125 ();
 sg13g2_decap_4 FILLER_30_132 ();
 sg13g2_fill_2 FILLER_30_136 ();
 sg13g2_fill_2 FILLER_30_156 ();
 sg13g2_fill_1 FILLER_30_158 ();
 sg13g2_decap_4 FILLER_30_164 ();
 sg13g2_fill_2 FILLER_30_188 ();
 sg13g2_decap_4 FILLER_30_193 ();
 sg13g2_fill_2 FILLER_30_197 ();
 sg13g2_decap_4 FILLER_30_203 ();
 sg13g2_fill_1 FILLER_30_207 ();
 sg13g2_fill_1 FILLER_30_230 ();
 sg13g2_fill_1 FILLER_30_241 ();
 sg13g2_fill_2 FILLER_30_252 ();
 sg13g2_fill_1 FILLER_30_254 ();
 sg13g2_fill_1 FILLER_30_267 ();
 sg13g2_fill_2 FILLER_30_296 ();
 sg13g2_fill_1 FILLER_30_303 ();
 sg13g2_fill_2 FILLER_30_314 ();
 sg13g2_fill_2 FILLER_30_321 ();
 sg13g2_fill_1 FILLER_30_323 ();
 sg13g2_fill_2 FILLER_30_328 ();
 sg13g2_fill_1 FILLER_30_330 ();
 sg13g2_fill_2 FILLER_30_389 ();
 sg13g2_fill_1 FILLER_30_391 ();
 sg13g2_fill_1 FILLER_30_410 ();
 sg13g2_fill_2 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_30_435 ();
 sg13g2_fill_1 FILLER_30_442 ();
 sg13g2_fill_2 FILLER_30_456 ();
 sg13g2_fill_2 FILLER_30_473 ();
 sg13g2_fill_1 FILLER_30_475 ();
 sg13g2_decap_8 FILLER_30_481 ();
 sg13g2_fill_1 FILLER_30_491 ();
 sg13g2_decap_8 FILLER_30_505 ();
 sg13g2_decap_4 FILLER_30_512 ();
 sg13g2_decap_4 FILLER_30_560 ();
 sg13g2_decap_8 FILLER_30_582 ();
 sg13g2_fill_2 FILLER_30_589 ();
 sg13g2_decap_8 FILLER_30_609 ();
 sg13g2_decap_4 FILLER_30_616 ();
 sg13g2_fill_1 FILLER_30_658 ();
 sg13g2_fill_2 FILLER_30_730 ();
 sg13g2_fill_2 FILLER_30_737 ();
 sg13g2_fill_1 FILLER_30_739 ();
 sg13g2_decap_4 FILLER_30_744 ();
 sg13g2_decap_8 FILLER_30_761 ();
 sg13g2_decap_8 FILLER_30_768 ();
 sg13g2_decap_4 FILLER_30_775 ();
 sg13g2_decap_8 FILLER_30_801 ();
 sg13g2_decap_8 FILLER_30_808 ();
 sg13g2_decap_4 FILLER_30_815 ();
 sg13g2_fill_1 FILLER_30_819 ();
 sg13g2_decap_4 FILLER_30_855 ();
 sg13g2_fill_2 FILLER_30_859 ();
 sg13g2_fill_1 FILLER_30_874 ();
 sg13g2_fill_2 FILLER_30_893 ();
 sg13g2_fill_1 FILLER_30_895 ();
 sg13g2_fill_2 FILLER_30_909 ();
 sg13g2_fill_1 FILLER_30_911 ();
 sg13g2_fill_1 FILLER_30_947 ();
 sg13g2_fill_2 FILLER_30_951 ();
 sg13g2_decap_8 FILLER_30_981 ();
 sg13g2_decap_8 FILLER_30_988 ();
 sg13g2_decap_8 FILLER_30_995 ();
 sg13g2_decap_8 FILLER_30_1002 ();
 sg13g2_decap_8 FILLER_30_1009 ();
 sg13g2_decap_8 FILLER_30_1016 ();
 sg13g2_decap_4 FILLER_30_1023 ();
 sg13g2_fill_2 FILLER_30_1027 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_4 ();
 sg13g2_fill_1 FILLER_31_32 ();
 sg13g2_decap_8 FILLER_31_50 ();
 sg13g2_decap_8 FILLER_31_57 ();
 sg13g2_decap_8 FILLER_31_64 ();
 sg13g2_fill_1 FILLER_31_71 ();
 sg13g2_fill_2 FILLER_31_82 ();
 sg13g2_fill_1 FILLER_31_84 ();
 sg13g2_fill_1 FILLER_31_94 ();
 sg13g2_fill_2 FILLER_31_100 ();
 sg13g2_decap_4 FILLER_31_137 ();
 sg13g2_fill_1 FILLER_31_141 ();
 sg13g2_fill_2 FILLER_31_211 ();
 sg13g2_fill_1 FILLER_31_213 ();
 sg13g2_fill_1 FILLER_31_228 ();
 sg13g2_decap_4 FILLER_31_238 ();
 sg13g2_fill_2 FILLER_31_242 ();
 sg13g2_decap_8 FILLER_31_264 ();
 sg13g2_decap_8 FILLER_31_271 ();
 sg13g2_fill_1 FILLER_31_278 ();
 sg13g2_fill_1 FILLER_31_284 ();
 sg13g2_decap_4 FILLER_31_298 ();
 sg13g2_fill_1 FILLER_31_302 ();
 sg13g2_fill_2 FILLER_31_313 ();
 sg13g2_decap_8 FILLER_31_325 ();
 sg13g2_decap_4 FILLER_31_332 ();
 sg13g2_fill_1 FILLER_31_336 ();
 sg13g2_fill_2 FILLER_31_342 ();
 sg13g2_fill_1 FILLER_31_347 ();
 sg13g2_fill_2 FILLER_31_376 ();
 sg13g2_fill_1 FILLER_31_391 ();
 sg13g2_decap_4 FILLER_31_421 ();
 sg13g2_fill_1 FILLER_31_425 ();
 sg13g2_decap_4 FILLER_31_454 ();
 sg13g2_fill_1 FILLER_31_458 ();
 sg13g2_fill_2 FILLER_31_469 ();
 sg13g2_decap_4 FILLER_31_486 ();
 sg13g2_fill_2 FILLER_31_490 ();
 sg13g2_decap_4 FILLER_31_520 ();
 sg13g2_fill_2 FILLER_31_528 ();
 sg13g2_fill_2 FILLER_31_560 ();
 sg13g2_decap_8 FILLER_31_589 ();
 sg13g2_fill_1 FILLER_31_596 ();
 sg13g2_fill_2 FILLER_31_611 ();
 sg13g2_fill_1 FILLER_31_613 ();
 sg13g2_fill_2 FILLER_31_619 ();
 sg13g2_decap_8 FILLER_31_626 ();
 sg13g2_fill_2 FILLER_31_633 ();
 sg13g2_decap_8 FILLER_31_648 ();
 sg13g2_decap_4 FILLER_31_655 ();
 sg13g2_fill_1 FILLER_31_659 ();
 sg13g2_decap_8 FILLER_31_664 ();
 sg13g2_fill_1 FILLER_31_671 ();
 sg13g2_fill_1 FILLER_31_686 ();
 sg13g2_fill_2 FILLER_31_696 ();
 sg13g2_fill_1 FILLER_31_708 ();
 sg13g2_fill_1 FILLER_31_718 ();
 sg13g2_decap_8 FILLER_31_732 ();
 sg13g2_decap_8 FILLER_31_739 ();
 sg13g2_fill_2 FILLER_31_746 ();
 sg13g2_decap_4 FILLER_31_772 ();
 sg13g2_fill_1 FILLER_31_776 ();
 sg13g2_fill_2 FILLER_31_790 ();
 sg13g2_fill_1 FILLER_31_792 ();
 sg13g2_decap_8 FILLER_31_803 ();
 sg13g2_fill_2 FILLER_31_810 ();
 sg13g2_fill_1 FILLER_31_827 ();
 sg13g2_fill_2 FILLER_31_832 ();
 sg13g2_fill_2 FILLER_31_843 ();
 sg13g2_fill_2 FILLER_31_923 ();
 sg13g2_decap_8 FILLER_31_935 ();
 sg13g2_decap_4 FILLER_31_942 ();
 sg13g2_fill_1 FILLER_31_946 ();
 sg13g2_decap_8 FILLER_31_950 ();
 sg13g2_decap_8 FILLER_31_957 ();
 sg13g2_decap_8 FILLER_31_964 ();
 sg13g2_decap_8 FILLER_31_971 ();
 sg13g2_decap_8 FILLER_31_978 ();
 sg13g2_decap_8 FILLER_31_985 ();
 sg13g2_decap_8 FILLER_31_992 ();
 sg13g2_decap_8 FILLER_31_999 ();
 sg13g2_decap_8 FILLER_31_1006 ();
 sg13g2_decap_8 FILLER_31_1013 ();
 sg13g2_decap_8 FILLER_31_1020 ();
 sg13g2_fill_2 FILLER_31_1027 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_7 ();
 sg13g2_decap_4 FILLER_32_15 ();
 sg13g2_fill_2 FILLER_32_19 ();
 sg13g2_decap_8 FILLER_32_62 ();
 sg13g2_fill_1 FILLER_32_69 ();
 sg13g2_decap_8 FILLER_32_79 ();
 sg13g2_decap_8 FILLER_32_86 ();
 sg13g2_decap_4 FILLER_32_93 ();
 sg13g2_fill_1 FILLER_32_97 ();
 sg13g2_fill_1 FILLER_32_115 ();
 sg13g2_decap_8 FILLER_32_125 ();
 sg13g2_fill_1 FILLER_32_132 ();
 sg13g2_fill_2 FILLER_32_148 ();
 sg13g2_decap_8 FILLER_32_164 ();
 sg13g2_decap_4 FILLER_32_171 ();
 sg13g2_decap_4 FILLER_32_188 ();
 sg13g2_fill_2 FILLER_32_192 ();
 sg13g2_fill_2 FILLER_32_222 ();
 sg13g2_decap_8 FILLER_32_229 ();
 sg13g2_fill_1 FILLER_32_236 ();
 sg13g2_decap_4 FILLER_32_266 ();
 sg13g2_decap_4 FILLER_32_345 ();
 sg13g2_fill_1 FILLER_32_349 ();
 sg13g2_decap_8 FILLER_32_376 ();
 sg13g2_fill_2 FILLER_32_383 ();
 sg13g2_fill_1 FILLER_32_385 ();
 sg13g2_fill_1 FILLER_32_406 ();
 sg13g2_decap_8 FILLER_32_412 ();
 sg13g2_decap_8 FILLER_32_419 ();
 sg13g2_fill_2 FILLER_32_426 ();
 sg13g2_fill_1 FILLER_32_428 ();
 sg13g2_decap_4 FILLER_32_451 ();
 sg13g2_fill_2 FILLER_32_455 ();
 sg13g2_decap_8 FILLER_32_476 ();
 sg13g2_decap_8 FILLER_32_483 ();
 sg13g2_decap_8 FILLER_32_490 ();
 sg13g2_fill_1 FILLER_32_510 ();
 sg13g2_fill_2 FILLER_32_515 ();
 sg13g2_fill_2 FILLER_32_530 ();
 sg13g2_fill_1 FILLER_32_562 ();
 sg13g2_decap_8 FILLER_32_583 ();
 sg13g2_fill_1 FILLER_32_590 ();
 sg13g2_fill_1 FILLER_32_605 ();
 sg13g2_decap_8 FILLER_32_647 ();
 sg13g2_fill_1 FILLER_32_654 ();
 sg13g2_fill_1 FILLER_32_668 ();
 sg13g2_fill_1 FILLER_32_682 ();
 sg13g2_decap_8 FILLER_32_721 ();
 sg13g2_fill_1 FILLER_32_741 ();
 sg13g2_fill_2 FILLER_32_767 ();
 sg13g2_fill_1 FILLER_32_800 ();
 sg13g2_decap_8 FILLER_32_826 ();
 sg13g2_decap_4 FILLER_32_833 ();
 sg13g2_fill_1 FILLER_32_837 ();
 sg13g2_decap_4 FILLER_32_843 ();
 sg13g2_decap_8 FILLER_32_854 ();
 sg13g2_decap_8 FILLER_32_861 ();
 sg13g2_fill_2 FILLER_32_868 ();
 sg13g2_fill_1 FILLER_32_896 ();
 sg13g2_fill_2 FILLER_32_905 ();
 sg13g2_decap_8 FILLER_32_920 ();
 sg13g2_decap_4 FILLER_32_931 ();
 sg13g2_decap_8 FILLER_32_961 ();
 sg13g2_decap_8 FILLER_32_968 ();
 sg13g2_decap_8 FILLER_32_975 ();
 sg13g2_decap_8 FILLER_32_982 ();
 sg13g2_decap_8 FILLER_32_989 ();
 sg13g2_decap_8 FILLER_32_996 ();
 sg13g2_decap_8 FILLER_32_1003 ();
 sg13g2_decap_8 FILLER_32_1010 ();
 sg13g2_decap_8 FILLER_32_1017 ();
 sg13g2_decap_4 FILLER_32_1024 ();
 sg13g2_fill_1 FILLER_32_1028 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_4 ();
 sg13g2_fill_2 FILLER_33_33 ();
 sg13g2_fill_2 FILLER_33_48 ();
 sg13g2_fill_1 FILLER_33_88 ();
 sg13g2_decap_4 FILLER_33_120 ();
 sg13g2_fill_1 FILLER_33_124 ();
 sg13g2_fill_2 FILLER_33_138 ();
 sg13g2_decap_8 FILLER_33_195 ();
 sg13g2_decap_8 FILLER_33_202 ();
 sg13g2_decap_4 FILLER_33_209 ();
 sg13g2_decap_4 FILLER_33_241 ();
 sg13g2_fill_1 FILLER_33_245 ();
 sg13g2_fill_2 FILLER_33_261 ();
 sg13g2_fill_1 FILLER_33_275 ();
 sg13g2_decap_8 FILLER_33_280 ();
 sg13g2_fill_2 FILLER_33_287 ();
 sg13g2_decap_4 FILLER_33_298 ();
 sg13g2_fill_2 FILLER_33_302 ();
 sg13g2_decap_8 FILLER_33_323 ();
 sg13g2_fill_1 FILLER_33_330 ();
 sg13g2_fill_2 FILLER_33_360 ();
 sg13g2_decap_4 FILLER_33_388 ();
 sg13g2_fill_1 FILLER_33_402 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_33_414 ();
 sg13g2_decap_4 FILLER_33_421 ();
 sg13g2_decap_4 FILLER_33_438 ();
 sg13g2_fill_1 FILLER_33_442 ();
 sg13g2_fill_2 FILLER_33_466 ();
 sg13g2_fill_2 FILLER_33_478 ();
 sg13g2_decap_4 FILLER_33_490 ();
 sg13g2_fill_2 FILLER_33_499 ();
 sg13g2_fill_2 FILLER_33_504 ();
 sg13g2_decap_8 FILLER_33_537 ();
 sg13g2_decap_8 FILLER_33_544 ();
 sg13g2_fill_1 FILLER_33_551 ();
 sg13g2_fill_2 FILLER_33_556 ();
 sg13g2_decap_4 FILLER_33_566 ();
 sg13g2_fill_2 FILLER_33_570 ();
 sg13g2_fill_1 FILLER_33_603 ();
 sg13g2_fill_1 FILLER_33_614 ();
 sg13g2_fill_1 FILLER_33_625 ();
 sg13g2_fill_2 FILLER_33_630 ();
 sg13g2_fill_2 FILLER_33_645 ();
 sg13g2_fill_1 FILLER_33_647 ();
 sg13g2_decap_8 FILLER_33_661 ();
 sg13g2_decap_8 FILLER_33_668 ();
 sg13g2_fill_2 FILLER_33_688 ();
 sg13g2_fill_1 FILLER_33_690 ();
 sg13g2_decap_4 FILLER_33_719 ();
 sg13g2_fill_1 FILLER_33_723 ();
 sg13g2_fill_2 FILLER_33_750 ();
 sg13g2_fill_1 FILLER_33_793 ();
 sg13g2_fill_1 FILLER_33_807 ();
 sg13g2_decap_8 FILLER_33_833 ();
 sg13g2_fill_1 FILLER_33_840 ();
 sg13g2_decap_4 FILLER_33_863 ();
 sg13g2_fill_1 FILLER_33_867 ();
 sg13g2_decap_4 FILLER_33_900 ();
 sg13g2_decap_8 FILLER_33_909 ();
 sg13g2_decap_4 FILLER_33_916 ();
 sg13g2_fill_2 FILLER_33_920 ();
 sg13g2_decap_8 FILLER_33_962 ();
 sg13g2_decap_8 FILLER_33_969 ();
 sg13g2_decap_8 FILLER_33_976 ();
 sg13g2_decap_8 FILLER_33_983 ();
 sg13g2_decap_8 FILLER_33_990 ();
 sg13g2_decap_8 FILLER_33_997 ();
 sg13g2_decap_8 FILLER_33_1004 ();
 sg13g2_decap_8 FILLER_33_1011 ();
 sg13g2_decap_8 FILLER_33_1018 ();
 sg13g2_decap_4 FILLER_33_1025 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_17 ();
 sg13g2_decap_4 FILLER_34_24 ();
 sg13g2_fill_2 FILLER_34_41 ();
 sg13g2_fill_1 FILLER_34_48 ();
 sg13g2_fill_2 FILLER_34_58 ();
 sg13g2_decap_8 FILLER_34_65 ();
 sg13g2_decap_8 FILLER_34_114 ();
 sg13g2_decap_4 FILLER_34_121 ();
 sg13g2_fill_1 FILLER_34_125 ();
 sg13g2_decap_8 FILLER_34_144 ();
 sg13g2_decap_4 FILLER_34_151 ();
 sg13g2_decap_8 FILLER_34_159 ();
 sg13g2_fill_2 FILLER_34_166 ();
 sg13g2_fill_1 FILLER_34_198 ();
 sg13g2_decap_4 FILLER_34_249 ();
 sg13g2_decap_8 FILLER_34_256 ();
 sg13g2_fill_1 FILLER_34_263 ();
 sg13g2_decap_8 FILLER_34_277 ();
 sg13g2_fill_2 FILLER_34_284 ();
 sg13g2_decap_8 FILLER_34_290 ();
 sg13g2_fill_2 FILLER_34_297 ();
 sg13g2_fill_1 FILLER_34_299 ();
 sg13g2_fill_2 FILLER_34_315 ();
 sg13g2_fill_1 FILLER_34_322 ();
 sg13g2_fill_1 FILLER_34_328 ();
 sg13g2_fill_2 FILLER_34_334 ();
 sg13g2_decap_8 FILLER_34_373 ();
 sg13g2_fill_2 FILLER_34_380 ();
 sg13g2_fill_1 FILLER_34_382 ();
 sg13g2_fill_2 FILLER_34_388 ();
 sg13g2_fill_1 FILLER_34_400 ();
 sg13g2_fill_1 FILLER_34_411 ();
 sg13g2_decap_4 FILLER_34_452 ();
 sg13g2_decap_8 FILLER_34_501 ();
 sg13g2_decap_4 FILLER_34_508 ();
 sg13g2_fill_2 FILLER_34_512 ();
 sg13g2_fill_1 FILLER_34_523 ();
 sg13g2_fill_2 FILLER_34_568 ();
 sg13g2_decap_4 FILLER_34_575 ();
 sg13g2_fill_1 FILLER_34_579 ();
 sg13g2_decap_8 FILLER_34_584 ();
 sg13g2_decap_8 FILLER_34_591 ();
 sg13g2_decap_8 FILLER_34_598 ();
 sg13g2_decap_8 FILLER_34_605 ();
 sg13g2_decap_8 FILLER_34_612 ();
 sg13g2_fill_1 FILLER_34_619 ();
 sg13g2_decap_4 FILLER_34_653 ();
 sg13g2_fill_1 FILLER_34_657 ();
 sg13g2_fill_2 FILLER_34_671 ();
 sg13g2_fill_1 FILLER_34_673 ();
 sg13g2_fill_2 FILLER_34_687 ();
 sg13g2_fill_1 FILLER_34_689 ();
 sg13g2_fill_2 FILLER_34_695 ();
 sg13g2_fill_1 FILLER_34_702 ();
 sg13g2_decap_8 FILLER_34_707 ();
 sg13g2_fill_1 FILLER_34_714 ();
 sg13g2_fill_2 FILLER_34_747 ();
 sg13g2_fill_2 FILLER_34_775 ();
 sg13g2_decap_4 FILLER_34_805 ();
 sg13g2_fill_1 FILLER_34_809 ();
 sg13g2_fill_2 FILLER_34_820 ();
 sg13g2_fill_1 FILLER_34_822 ();
 sg13g2_decap_8 FILLER_34_837 ();
 sg13g2_decap_8 FILLER_34_894 ();
 sg13g2_fill_2 FILLER_34_906 ();
 sg13g2_fill_1 FILLER_34_908 ();
 sg13g2_decap_8 FILLER_34_935 ();
 sg13g2_decap_8 FILLER_34_942 ();
 sg13g2_decap_8 FILLER_34_949 ();
 sg13g2_decap_8 FILLER_34_956 ();
 sg13g2_decap_8 FILLER_34_963 ();
 sg13g2_decap_8 FILLER_34_970 ();
 sg13g2_decap_8 FILLER_34_977 ();
 sg13g2_decap_8 FILLER_34_984 ();
 sg13g2_decap_8 FILLER_34_991 ();
 sg13g2_decap_8 FILLER_34_998 ();
 sg13g2_decap_8 FILLER_34_1005 ();
 sg13g2_decap_8 FILLER_34_1012 ();
 sg13g2_decap_8 FILLER_34_1019 ();
 sg13g2_fill_2 FILLER_34_1026 ();
 sg13g2_fill_1 FILLER_34_1028 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_7 ();
 sg13g2_decap_4 FILLER_35_62 ();
 sg13g2_decap_4 FILLER_35_71 ();
 sg13g2_fill_1 FILLER_35_75 ();
 sg13g2_decap_4 FILLER_35_86 ();
 sg13g2_fill_1 FILLER_35_90 ();
 sg13g2_decap_8 FILLER_35_96 ();
 sg13g2_fill_2 FILLER_35_103 ();
 sg13g2_decap_4 FILLER_35_133 ();
 sg13g2_fill_2 FILLER_35_137 ();
 sg13g2_fill_2 FILLER_35_154 ();
 sg13g2_fill_2 FILLER_35_165 ();
 sg13g2_fill_1 FILLER_35_167 ();
 sg13g2_fill_2 FILLER_35_171 ();
 sg13g2_decap_8 FILLER_35_214 ();
 sg13g2_fill_1 FILLER_35_221 ();
 sg13g2_decap_8 FILLER_35_251 ();
 sg13g2_fill_1 FILLER_35_258 ();
 sg13g2_fill_2 FILLER_35_324 ();
 sg13g2_fill_1 FILLER_35_339 ();
 sg13g2_decap_8 FILLER_35_360 ();
 sg13g2_decap_4 FILLER_35_393 ();
 sg13g2_fill_1 FILLER_35_402 ();
 sg13g2_decap_8 FILLER_35_418 ();
 sg13g2_decap_8 FILLER_35_425 ();
 sg13g2_decap_4 FILLER_35_432 ();
 sg13g2_fill_2 FILLER_35_436 ();
 sg13g2_decap_8 FILLER_35_456 ();
 sg13g2_decap_8 FILLER_35_463 ();
 sg13g2_decap_8 FILLER_35_470 ();
 sg13g2_fill_2 FILLER_35_477 ();
 sg13g2_decap_8 FILLER_35_494 ();
 sg13g2_fill_2 FILLER_35_501 ();
 sg13g2_decap_8 FILLER_35_507 ();
 sg13g2_fill_2 FILLER_35_514 ();
 sg13g2_fill_1 FILLER_35_546 ();
 sg13g2_fill_2 FILLER_35_561 ();
 sg13g2_fill_1 FILLER_35_563 ();
 sg13g2_decap_8 FILLER_35_581 ();
 sg13g2_decap_8 FILLER_35_588 ();
 sg13g2_decap_8 FILLER_35_595 ();
 sg13g2_fill_2 FILLER_35_602 ();
 sg13g2_fill_2 FILLER_35_617 ();
 sg13g2_fill_2 FILLER_35_632 ();
 sg13g2_fill_1 FILLER_35_634 ();
 sg13g2_fill_2 FILLER_35_644 ();
 sg13g2_fill_1 FILLER_35_646 ();
 sg13g2_fill_2 FILLER_35_670 ();
 sg13g2_decap_8 FILLER_35_689 ();
 sg13g2_decap_4 FILLER_35_696 ();
 sg13g2_fill_2 FILLER_35_700 ();
 sg13g2_decap_4 FILLER_35_715 ();
 sg13g2_fill_1 FILLER_35_719 ();
 sg13g2_decap_8 FILLER_35_737 ();
 sg13g2_decap_8 FILLER_35_744 ();
 sg13g2_decap_4 FILLER_35_751 ();
 sg13g2_fill_2 FILLER_35_775 ();
 sg13g2_decap_4 FILLER_35_790 ();
 sg13g2_fill_2 FILLER_35_794 ();
 sg13g2_decap_8 FILLER_35_809 ();
 sg13g2_decap_8 FILLER_35_816 ();
 sg13g2_decap_8 FILLER_35_842 ();
 sg13g2_fill_2 FILLER_35_849 ();
 sg13g2_decap_8 FILLER_35_859 ();
 sg13g2_fill_2 FILLER_35_866 ();
 sg13g2_fill_1 FILLER_35_873 ();
 sg13g2_decap_8 FILLER_35_889 ();
 sg13g2_fill_1 FILLER_35_921 ();
 sg13g2_decap_8 FILLER_35_950 ();
 sg13g2_decap_8 FILLER_35_957 ();
 sg13g2_decap_8 FILLER_35_964 ();
 sg13g2_decap_8 FILLER_35_971 ();
 sg13g2_decap_8 FILLER_35_978 ();
 sg13g2_decap_8 FILLER_35_985 ();
 sg13g2_decap_8 FILLER_35_992 ();
 sg13g2_decap_8 FILLER_35_999 ();
 sg13g2_decap_8 FILLER_35_1006 ();
 sg13g2_decap_8 FILLER_35_1013 ();
 sg13g2_decap_8 FILLER_35_1020 ();
 sg13g2_fill_2 FILLER_35_1027 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_11 ();
 sg13g2_decap_8 FILLER_36_17 ();
 sg13g2_decap_4 FILLER_36_24 ();
 sg13g2_decap_8 FILLER_36_57 ();
 sg13g2_decap_4 FILLER_36_64 ();
 sg13g2_fill_2 FILLER_36_68 ();
 sg13g2_fill_2 FILLER_36_93 ();
 sg13g2_fill_1 FILLER_36_95 ();
 sg13g2_fill_2 FILLER_36_104 ();
 sg13g2_fill_1 FILLER_36_106 ();
 sg13g2_decap_4 FILLER_36_133 ();
 sg13g2_fill_1 FILLER_36_137 ();
 sg13g2_fill_2 FILLER_36_158 ();
 sg13g2_fill_1 FILLER_36_160 ();
 sg13g2_decap_4 FILLER_36_171 ();
 sg13g2_fill_2 FILLER_36_175 ();
 sg13g2_fill_2 FILLER_36_190 ();
 sg13g2_fill_1 FILLER_36_192 ();
 sg13g2_fill_1 FILLER_36_197 ();
 sg13g2_fill_2 FILLER_36_278 ();
 sg13g2_decap_8 FILLER_36_310 ();
 sg13g2_decap_4 FILLER_36_317 ();
 sg13g2_fill_2 FILLER_36_321 ();
 sg13g2_decap_8 FILLER_36_338 ();
 sg13g2_decap_8 FILLER_36_372 ();
 sg13g2_decap_4 FILLER_36_379 ();
 sg13g2_fill_2 FILLER_36_396 ();
 sg13g2_decap_4 FILLER_36_418 ();
 sg13g2_fill_2 FILLER_36_422 ();
 sg13g2_decap_8 FILLER_36_428 ();
 sg13g2_decap_8 FILLER_36_435 ();
 sg13g2_decap_8 FILLER_36_442 ();
 sg13g2_fill_2 FILLER_36_449 ();
 sg13g2_fill_1 FILLER_36_451 ();
 sg13g2_decap_8 FILLER_36_456 ();
 sg13g2_fill_2 FILLER_36_463 ();
 sg13g2_fill_1 FILLER_36_497 ();
 sg13g2_decap_8 FILLER_36_525 ();
 sg13g2_decap_8 FILLER_36_532 ();
 sg13g2_fill_1 FILLER_36_539 ();
 sg13g2_fill_2 FILLER_36_569 ();
 sg13g2_decap_4 FILLER_36_581 ();
 sg13g2_decap_8 FILLER_36_628 ();
 sg13g2_fill_1 FILLER_36_635 ();
 sg13g2_fill_2 FILLER_36_666 ();
 sg13g2_decap_8 FILLER_36_716 ();
 sg13g2_decap_4 FILLER_36_755 ();
 sg13g2_decap_4 FILLER_36_785 ();
 sg13g2_fill_1 FILLER_36_789 ();
 sg13g2_decap_8 FILLER_36_801 ();
 sg13g2_decap_8 FILLER_36_808 ();
 sg13g2_fill_1 FILLER_36_834 ();
 sg13g2_decap_8 FILLER_36_848 ();
 sg13g2_decap_4 FILLER_36_855 ();
 sg13g2_fill_2 FILLER_36_859 ();
 sg13g2_fill_1 FILLER_36_907 ();
 sg13g2_decap_8 FILLER_36_945 ();
 sg13g2_decap_8 FILLER_36_952 ();
 sg13g2_decap_8 FILLER_36_959 ();
 sg13g2_decap_8 FILLER_36_966 ();
 sg13g2_decap_8 FILLER_36_973 ();
 sg13g2_decap_8 FILLER_36_980 ();
 sg13g2_decap_8 FILLER_36_987 ();
 sg13g2_decap_8 FILLER_36_994 ();
 sg13g2_decap_8 FILLER_36_1001 ();
 sg13g2_decap_8 FILLER_36_1008 ();
 sg13g2_decap_8 FILLER_36_1015 ();
 sg13g2_decap_8 FILLER_36_1022 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_decap_4 FILLER_37_32 ();
 sg13g2_fill_2 FILLER_37_36 ();
 sg13g2_fill_1 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_55 ();
 sg13g2_decap_8 FILLER_37_62 ();
 sg13g2_fill_2 FILLER_37_69 ();
 sg13g2_decap_8 FILLER_37_95 ();
 sg13g2_fill_2 FILLER_37_102 ();
 sg13g2_fill_1 FILLER_37_104 ();
 sg13g2_decap_4 FILLER_37_118 ();
 sg13g2_fill_2 FILLER_37_122 ();
 sg13g2_decap_8 FILLER_37_137 ();
 sg13g2_fill_2 FILLER_37_144 ();
 sg13g2_fill_2 FILLER_37_164 ();
 sg13g2_fill_1 FILLER_37_166 ();
 sg13g2_decap_8 FILLER_37_170 ();
 sg13g2_decap_8 FILLER_37_177 ();
 sg13g2_decap_8 FILLER_37_184 ();
 sg13g2_decap_8 FILLER_37_191 ();
 sg13g2_decap_4 FILLER_37_198 ();
 sg13g2_fill_1 FILLER_37_202 ();
 sg13g2_decap_8 FILLER_37_207 ();
 sg13g2_decap_8 FILLER_37_214 ();
 sg13g2_decap_8 FILLER_37_221 ();
 sg13g2_decap_8 FILLER_37_228 ();
 sg13g2_decap_8 FILLER_37_235 ();
 sg13g2_fill_2 FILLER_37_242 ();
 sg13g2_fill_1 FILLER_37_244 ();
 sg13g2_decap_8 FILLER_37_260 ();
 sg13g2_fill_2 FILLER_37_267 ();
 sg13g2_fill_2 FILLER_37_309 ();
 sg13g2_fill_1 FILLER_37_311 ();
 sg13g2_fill_2 FILLER_37_317 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_fill_2 FILLER_37_364 ();
 sg13g2_decap_4 FILLER_37_392 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_4 FILLER_37_414 ();
 sg13g2_fill_1 FILLER_37_418 ();
 sg13g2_fill_1 FILLER_37_446 ();
 sg13g2_decap_8 FILLER_37_493 ();
 sg13g2_decap_8 FILLER_37_500 ();
 sg13g2_decap_8 FILLER_37_507 ();
 sg13g2_decap_4 FILLER_37_514 ();
 sg13g2_fill_2 FILLER_37_518 ();
 sg13g2_decap_4 FILLER_37_533 ();
 sg13g2_fill_1 FILLER_37_537 ();
 sg13g2_decap_8 FILLER_37_558 ();
 sg13g2_fill_2 FILLER_37_565 ();
 sg13g2_fill_1 FILLER_37_567 ();
 sg13g2_decap_4 FILLER_37_572 ();
 sg13g2_fill_2 FILLER_37_576 ();
 sg13g2_decap_4 FILLER_37_631 ();
 sg13g2_fill_1 FILLER_37_635 ();
 sg13g2_fill_2 FILLER_37_645 ();
 sg13g2_fill_2 FILLER_37_657 ();
 sg13g2_fill_2 FILLER_37_664 ();
 sg13g2_fill_1 FILLER_37_666 ();
 sg13g2_fill_1 FILLER_37_672 ();
 sg13g2_fill_1 FILLER_37_679 ();
 sg13g2_decap_4 FILLER_37_697 ();
 sg13g2_decap_8 FILLER_37_718 ();
 sg13g2_fill_2 FILLER_37_725 ();
 sg13g2_decap_4 FILLER_37_743 ();
 sg13g2_fill_1 FILLER_37_747 ();
 sg13g2_decap_8 FILLER_37_782 ();
 sg13g2_fill_2 FILLER_37_808 ();
 sg13g2_decap_8 FILLER_37_814 ();
 sg13g2_fill_1 FILLER_37_821 ();
 sg13g2_decap_4 FILLER_37_839 ();
 sg13g2_fill_1 FILLER_37_843 ();
 sg13g2_decap_8 FILLER_37_849 ();
 sg13g2_decap_8 FILLER_37_856 ();
 sg13g2_fill_2 FILLER_37_863 ();
 sg13g2_fill_1 FILLER_37_865 ();
 sg13g2_fill_1 FILLER_37_881 ();
 sg13g2_fill_2 FILLER_37_890 ();
 sg13g2_fill_1 FILLER_37_892 ();
 sg13g2_fill_1 FILLER_37_921 ();
 sg13g2_fill_1 FILLER_37_926 ();
 sg13g2_decap_8 FILLER_37_936 ();
 sg13g2_decap_8 FILLER_37_943 ();
 sg13g2_decap_8 FILLER_37_950 ();
 sg13g2_decap_8 FILLER_37_957 ();
 sg13g2_decap_8 FILLER_37_964 ();
 sg13g2_decap_8 FILLER_37_971 ();
 sg13g2_decap_8 FILLER_37_978 ();
 sg13g2_decap_8 FILLER_37_985 ();
 sg13g2_decap_8 FILLER_37_992 ();
 sg13g2_decap_8 FILLER_37_999 ();
 sg13g2_decap_8 FILLER_37_1006 ();
 sg13g2_decap_8 FILLER_37_1013 ();
 sg13g2_decap_8 FILLER_37_1020 ();
 sg13g2_fill_2 FILLER_37_1027 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_13 ();
 sg13g2_fill_2 FILLER_38_20 ();
 sg13g2_fill_2 FILLER_38_40 ();
 sg13g2_fill_1 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_60 ();
 sg13g2_decap_8 FILLER_38_92 ();
 sg13g2_fill_1 FILLER_38_99 ();
 sg13g2_fill_2 FILLER_38_121 ();
 sg13g2_fill_1 FILLER_38_123 ();
 sg13g2_decap_4 FILLER_38_150 ();
 sg13g2_fill_1 FILLER_38_154 ();
 sg13g2_fill_2 FILLER_38_166 ();
 sg13g2_fill_1 FILLER_38_173 ();
 sg13g2_fill_1 FILLER_38_179 ();
 sg13g2_decap_4 FILLER_38_185 ();
 sg13g2_fill_2 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_195 ();
 sg13g2_decap_4 FILLER_38_202 ();
 sg13g2_fill_1 FILLER_38_246 ();
 sg13g2_decap_4 FILLER_38_270 ();
 sg13g2_decap_8 FILLER_38_278 ();
 sg13g2_decap_8 FILLER_38_285 ();
 sg13g2_fill_2 FILLER_38_305 ();
 sg13g2_fill_1 FILLER_38_307 ();
 sg13g2_decap_4 FILLER_38_321 ();
 sg13g2_decap_4 FILLER_38_330 ();
 sg13g2_fill_2 FILLER_38_334 ();
 sg13g2_fill_1 FILLER_38_376 ();
 sg13g2_fill_1 FILLER_38_390 ();
 sg13g2_fill_1 FILLER_38_397 ();
 sg13g2_fill_2 FILLER_38_403 ();
 sg13g2_fill_1 FILLER_38_405 ();
 sg13g2_fill_1 FILLER_38_420 ();
 sg13g2_decap_8 FILLER_38_461 ();
 sg13g2_decap_4 FILLER_38_468 ();
 sg13g2_fill_1 FILLER_38_476 ();
 sg13g2_fill_2 FILLER_38_482 ();
 sg13g2_fill_1 FILLER_38_493 ();
 sg13g2_fill_2 FILLER_38_566 ();
 sg13g2_fill_1 FILLER_38_572 ();
 sg13g2_fill_1 FILLER_38_582 ();
 sg13g2_fill_2 FILLER_38_586 ();
 sg13g2_fill_1 FILLER_38_592 ();
 sg13g2_fill_1 FILLER_38_621 ();
 sg13g2_decap_8 FILLER_38_659 ();
 sg13g2_fill_1 FILLER_38_676 ();
 sg13g2_decap_4 FILLER_38_690 ();
 sg13g2_fill_1 FILLER_38_709 ();
 sg13g2_fill_2 FILLER_38_713 ();
 sg13g2_fill_1 FILLER_38_715 ();
 sg13g2_decap_4 FILLER_38_725 ();
 sg13g2_fill_1 FILLER_38_729 ();
 sg13g2_decap_8 FILLER_38_739 ();
 sg13g2_fill_2 FILLER_38_746 ();
 sg13g2_fill_1 FILLER_38_748 ();
 sg13g2_decap_4 FILLER_38_778 ();
 sg13g2_decap_8 FILLER_38_787 ();
 sg13g2_fill_1 FILLER_38_794 ();
 sg13g2_fill_2 FILLER_38_803 ();
 sg13g2_decap_8 FILLER_38_825 ();
 sg13g2_decap_4 FILLER_38_832 ();
 sg13g2_decap_4 FILLER_38_841 ();
 sg13g2_fill_2 FILLER_38_850 ();
 sg13g2_fill_1 FILLER_38_852 ();
 sg13g2_fill_1 FILLER_38_882 ();
 sg13g2_fill_2 FILLER_38_897 ();
 sg13g2_fill_1 FILLER_38_899 ();
 sg13g2_fill_1 FILLER_38_914 ();
 sg13g2_decap_8 FILLER_38_919 ();
 sg13g2_decap_8 FILLER_38_926 ();
 sg13g2_decap_8 FILLER_38_933 ();
 sg13g2_decap_8 FILLER_38_940 ();
 sg13g2_decap_8 FILLER_38_947 ();
 sg13g2_decap_8 FILLER_38_954 ();
 sg13g2_decap_8 FILLER_38_961 ();
 sg13g2_decap_8 FILLER_38_968 ();
 sg13g2_decap_8 FILLER_38_975 ();
 sg13g2_decap_8 FILLER_38_982 ();
 sg13g2_decap_8 FILLER_38_989 ();
 sg13g2_decap_8 FILLER_38_996 ();
 sg13g2_decap_8 FILLER_38_1003 ();
 sg13g2_decap_8 FILLER_38_1010 ();
 sg13g2_decap_8 FILLER_38_1017 ();
 sg13g2_decap_4 FILLER_38_1024 ();
 sg13g2_fill_1 FILLER_38_1028 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_2 ();
 sg13g2_decap_4 FILLER_39_61 ();
 sg13g2_fill_2 FILLER_39_65 ();
 sg13g2_decap_8 FILLER_39_80 ();
 sg13g2_fill_1 FILLER_39_126 ();
 sg13g2_fill_2 FILLER_39_131 ();
 sg13g2_fill_2 FILLER_39_146 ();
 sg13g2_fill_2 FILLER_39_184 ();
 sg13g2_fill_2 FILLER_39_214 ();
 sg13g2_fill_2 FILLER_39_233 ();
 sg13g2_fill_2 FILLER_39_240 ();
 sg13g2_decap_4 FILLER_39_260 ();
 sg13g2_fill_1 FILLER_39_264 ();
 sg13g2_fill_2 FILLER_39_269 ();
 sg13g2_fill_1 FILLER_39_271 ();
 sg13g2_fill_2 FILLER_39_312 ();
 sg13g2_fill_1 FILLER_39_314 ();
 sg13g2_decap_8 FILLER_39_325 ();
 sg13g2_decap_4 FILLER_39_332 ();
 sg13g2_fill_1 FILLER_39_336 ();
 sg13g2_decap_8 FILLER_39_350 ();
 sg13g2_fill_1 FILLER_39_357 ();
 sg13g2_fill_1 FILLER_39_398 ();
 sg13g2_decap_8 FILLER_39_404 ();
 sg13g2_fill_1 FILLER_39_411 ();
 sg13g2_decap_8 FILLER_39_416 ();
 sg13g2_fill_2 FILLER_39_423 ();
 sg13g2_fill_1 FILLER_39_425 ();
 sg13g2_fill_2 FILLER_39_430 ();
 sg13g2_fill_2 FILLER_39_445 ();
 sg13g2_decap_4 FILLER_39_452 ();
 sg13g2_fill_2 FILLER_39_456 ();
 sg13g2_fill_1 FILLER_39_498 ();
 sg13g2_decap_8 FILLER_39_503 ();
 sg13g2_decap_8 FILLER_39_510 ();
 sg13g2_fill_1 FILLER_39_517 ();
 sg13g2_decap_8 FILLER_39_531 ();
 sg13g2_fill_1 FILLER_39_538 ();
 sg13g2_fill_2 FILLER_39_548 ();
 sg13g2_fill_1 FILLER_39_550 ();
 sg13g2_fill_1 FILLER_39_556 ();
 sg13g2_fill_1 FILLER_39_581 ();
 sg13g2_decap_8 FILLER_39_615 ();
 sg13g2_fill_1 FILLER_39_622 ();
 sg13g2_fill_1 FILLER_39_635 ();
 sg13g2_fill_1 FILLER_39_664 ();
 sg13g2_fill_2 FILLER_39_693 ();
 sg13g2_fill_2 FILLER_39_705 ();
 sg13g2_fill_1 FILLER_39_712 ();
 sg13g2_fill_1 FILLER_39_740 ();
 sg13g2_decap_8 FILLER_39_746 ();
 sg13g2_fill_2 FILLER_39_753 ();
 sg13g2_decap_4 FILLER_39_770 ();
 sg13g2_fill_2 FILLER_39_774 ();
 sg13g2_fill_1 FILLER_39_796 ();
 sg13g2_fill_2 FILLER_39_814 ();
 sg13g2_fill_1 FILLER_39_816 ();
 sg13g2_fill_2 FILLER_39_832 ();
 sg13g2_fill_2 FILLER_39_839 ();
 sg13g2_fill_1 FILLER_39_841 ();
 sg13g2_fill_2 FILLER_39_882 ();
 sg13g2_decap_4 FILLER_39_906 ();
 sg13g2_decap_8 FILLER_39_937 ();
 sg13g2_decap_8 FILLER_39_944 ();
 sg13g2_decap_8 FILLER_39_951 ();
 sg13g2_decap_8 FILLER_39_958 ();
 sg13g2_decap_8 FILLER_39_965 ();
 sg13g2_decap_8 FILLER_39_972 ();
 sg13g2_decap_8 FILLER_39_979 ();
 sg13g2_decap_8 FILLER_39_986 ();
 sg13g2_decap_8 FILLER_39_993 ();
 sg13g2_decap_8 FILLER_39_1000 ();
 sg13g2_decap_8 FILLER_39_1007 ();
 sg13g2_decap_8 FILLER_39_1014 ();
 sg13g2_decap_8 FILLER_39_1021 ();
 sg13g2_fill_1 FILLER_39_1028 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_12 ();
 sg13g2_decap_8 FILLER_40_19 ();
 sg13g2_decap_4 FILLER_40_26 ();
 sg13g2_fill_1 FILLER_40_30 ();
 sg13g2_decap_4 FILLER_40_35 ();
 sg13g2_fill_1 FILLER_40_39 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_4 FILLER_40_56 ();
 sg13g2_fill_1 FILLER_40_78 ();
 sg13g2_decap_8 FILLER_40_88 ();
 sg13g2_fill_2 FILLER_40_95 ();
 sg13g2_fill_2 FILLER_40_102 ();
 sg13g2_decap_8 FILLER_40_107 ();
 sg13g2_decap_8 FILLER_40_114 ();
 sg13g2_decap_8 FILLER_40_121 ();
 sg13g2_decap_8 FILLER_40_128 ();
 sg13g2_fill_2 FILLER_40_135 ();
 sg13g2_fill_2 FILLER_40_150 ();
 sg13g2_fill_1 FILLER_40_152 ();
 sg13g2_decap_8 FILLER_40_162 ();
 sg13g2_fill_2 FILLER_40_169 ();
 sg13g2_fill_1 FILLER_40_171 ();
 sg13g2_fill_1 FILLER_40_182 ();
 sg13g2_decap_8 FILLER_40_186 ();
 sg13g2_decap_8 FILLER_40_193 ();
 sg13g2_decap_8 FILLER_40_200 ();
 sg13g2_decap_8 FILLER_40_207 ();
 sg13g2_decap_8 FILLER_40_214 ();
 sg13g2_fill_2 FILLER_40_221 ();
 sg13g2_fill_1 FILLER_40_227 ();
 sg13g2_fill_1 FILLER_40_233 ();
 sg13g2_decap_8 FILLER_40_243 ();
 sg13g2_decap_8 FILLER_40_283 ();
 sg13g2_decap_8 FILLER_40_290 ();
 sg13g2_fill_1 FILLER_40_297 ();
 sg13g2_decap_4 FILLER_40_302 ();
 sg13g2_fill_2 FILLER_40_306 ();
 sg13g2_fill_2 FILLER_40_318 ();
 sg13g2_fill_2 FILLER_40_351 ();
 sg13g2_fill_1 FILLER_40_353 ();
 sg13g2_fill_2 FILLER_40_367 ();
 sg13g2_fill_1 FILLER_40_382 ();
 sg13g2_decap_8 FILLER_40_393 ();
 sg13g2_decap_8 FILLER_40_400 ();
 sg13g2_fill_2 FILLER_40_444 ();
 sg13g2_decap_8 FILLER_40_478 ();
 sg13g2_decap_4 FILLER_40_485 ();
 sg13g2_fill_1 FILLER_40_489 ();
 sg13g2_fill_1 FILLER_40_494 ();
 sg13g2_decap_8 FILLER_40_504 ();
 sg13g2_fill_1 FILLER_40_511 ();
 sg13g2_decap_8 FILLER_40_530 ();
 sg13g2_fill_2 FILLER_40_537 ();
 sg13g2_fill_2 FILLER_40_544 ();
 sg13g2_fill_1 FILLER_40_546 ();
 sg13g2_fill_2 FILLER_40_564 ();
 sg13g2_fill_1 FILLER_40_566 ();
 sg13g2_decap_8 FILLER_40_571 ();
 sg13g2_decap_8 FILLER_40_578 ();
 sg13g2_fill_2 FILLER_40_585 ();
 sg13g2_fill_2 FILLER_40_607 ();
 sg13g2_decap_8 FILLER_40_618 ();
 sg13g2_decap_4 FILLER_40_625 ();
 sg13g2_fill_2 FILLER_40_629 ();
 sg13g2_decap_8 FILLER_40_653 ();
 sg13g2_decap_4 FILLER_40_660 ();
 sg13g2_fill_2 FILLER_40_664 ();
 sg13g2_decap_8 FILLER_40_679 ();
 sg13g2_decap_8 FILLER_40_686 ();
 sg13g2_fill_2 FILLER_40_693 ();
 sg13g2_fill_2 FILLER_40_709 ();
 sg13g2_fill_1 FILLER_40_711 ();
 sg13g2_decap_8 FILLER_40_730 ();
 sg13g2_fill_2 FILLER_40_737 ();
 sg13g2_fill_1 FILLER_40_739 ();
 sg13g2_fill_2 FILLER_40_745 ();
 sg13g2_decap_4 FILLER_40_778 ();
 sg13g2_decap_8 FILLER_40_786 ();
 sg13g2_fill_1 FILLER_40_812 ();
 sg13g2_decap_4 FILLER_40_852 ();
 sg13g2_fill_1 FILLER_40_856 ();
 sg13g2_decap_4 FILLER_40_870 ();
 sg13g2_fill_2 FILLER_40_874 ();
 sg13g2_fill_2 FILLER_40_880 ();
 sg13g2_decap_8 FILLER_40_909 ();
 sg13g2_decap_4 FILLER_40_916 ();
 sg13g2_fill_2 FILLER_40_920 ();
 sg13g2_decap_8 FILLER_40_931 ();
 sg13g2_decap_8 FILLER_40_938 ();
 sg13g2_decap_8 FILLER_40_945 ();
 sg13g2_decap_8 FILLER_40_952 ();
 sg13g2_decap_8 FILLER_40_959 ();
 sg13g2_decap_8 FILLER_40_966 ();
 sg13g2_decap_8 FILLER_40_973 ();
 sg13g2_decap_8 FILLER_40_980 ();
 sg13g2_decap_8 FILLER_40_987 ();
 sg13g2_decap_8 FILLER_40_994 ();
 sg13g2_decap_8 FILLER_40_1001 ();
 sg13g2_decap_8 FILLER_40_1008 ();
 sg13g2_decap_8 FILLER_40_1015 ();
 sg13g2_decap_8 FILLER_40_1022 ();
 sg13g2_fill_2 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_2 ();
 sg13g2_fill_2 FILLER_41_36 ();
 sg13g2_decap_4 FILLER_41_50 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_fill_1 FILLER_41_91 ();
 sg13g2_decap_4 FILLER_41_114 ();
 sg13g2_fill_1 FILLER_41_118 ();
 sg13g2_fill_1 FILLER_41_145 ();
 sg13g2_fill_2 FILLER_41_156 ();
 sg13g2_fill_1 FILLER_41_158 ();
 sg13g2_decap_8 FILLER_41_169 ();
 sg13g2_fill_2 FILLER_41_181 ();
 sg13g2_fill_2 FILLER_41_223 ();
 sg13g2_fill_1 FILLER_41_225 ();
 sg13g2_fill_1 FILLER_41_240 ();
 sg13g2_fill_1 FILLER_41_250 ();
 sg13g2_fill_1 FILLER_41_278 ();
 sg13g2_fill_2 FILLER_41_292 ();
 sg13g2_fill_1 FILLER_41_294 ();
 sg13g2_fill_2 FILLER_41_327 ();
 sg13g2_decap_8 FILLER_41_338 ();
 sg13g2_decap_8 FILLER_41_345 ();
 sg13g2_decap_4 FILLER_41_352 ();
 sg13g2_fill_2 FILLER_41_374 ();
 sg13g2_decap_4 FILLER_41_391 ();
 sg13g2_fill_2 FILLER_41_408 ();
 sg13g2_fill_1 FILLER_41_410 ();
 sg13g2_fill_1 FILLER_41_415 ();
 sg13g2_fill_1 FILLER_41_429 ();
 sg13g2_decap_8 FILLER_41_439 ();
 sg13g2_decap_8 FILLER_41_446 ();
 sg13g2_fill_2 FILLER_41_453 ();
 sg13g2_fill_1 FILLER_41_455 ();
 sg13g2_decap_4 FILLER_41_477 ();
 sg13g2_fill_2 FILLER_41_481 ();
 sg13g2_decap_4 FILLER_41_510 ();
 sg13g2_fill_1 FILLER_41_527 ();
 sg13g2_decap_8 FILLER_41_570 ();
 sg13g2_fill_2 FILLER_41_577 ();
 sg13g2_decap_4 FILLER_41_599 ();
 sg13g2_decap_8 FILLER_41_620 ();
 sg13g2_decap_4 FILLER_41_627 ();
 sg13g2_decap_8 FILLER_41_656 ();
 sg13g2_fill_2 FILLER_41_663 ();
 sg13g2_decap_4 FILLER_41_681 ();
 sg13g2_fill_1 FILLER_41_685 ();
 sg13g2_decap_8 FILLER_41_718 ();
 sg13g2_decap_8 FILLER_41_725 ();
 sg13g2_fill_2 FILLER_41_732 ();
 sg13g2_fill_1 FILLER_41_734 ();
 sg13g2_fill_1 FILLER_41_762 ();
 sg13g2_decap_4 FILLER_41_782 ();
 sg13g2_fill_2 FILLER_41_786 ();
 sg13g2_decap_8 FILLER_41_815 ();
 sg13g2_decap_8 FILLER_41_822 ();
 sg13g2_decap_8 FILLER_41_829 ();
 sg13g2_decap_8 FILLER_41_836 ();
 sg13g2_decap_4 FILLER_41_843 ();
 sg13g2_fill_1 FILLER_41_847 ();
 sg13g2_decap_8 FILLER_41_876 ();
 sg13g2_decap_4 FILLER_41_883 ();
 sg13g2_decap_8 FILLER_41_891 ();
 sg13g2_decap_8 FILLER_41_898 ();
 sg13g2_decap_8 FILLER_41_905 ();
 sg13g2_decap_8 FILLER_41_912 ();
 sg13g2_decap_8 FILLER_41_919 ();
 sg13g2_decap_8 FILLER_41_926 ();
 sg13g2_decap_8 FILLER_41_933 ();
 sg13g2_decap_8 FILLER_41_940 ();
 sg13g2_decap_8 FILLER_41_947 ();
 sg13g2_decap_8 FILLER_41_954 ();
 sg13g2_decap_8 FILLER_41_961 ();
 sg13g2_decap_8 FILLER_41_968 ();
 sg13g2_decap_8 FILLER_41_975 ();
 sg13g2_decap_8 FILLER_41_982 ();
 sg13g2_decap_8 FILLER_41_989 ();
 sg13g2_decap_8 FILLER_41_996 ();
 sg13g2_decap_8 FILLER_41_1003 ();
 sg13g2_decap_8 FILLER_41_1010 ();
 sg13g2_decap_8 FILLER_41_1017 ();
 sg13g2_decap_4 FILLER_41_1024 ();
 sg13g2_fill_1 FILLER_41_1028 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_13 ();
 sg13g2_decap_4 FILLER_42_20 ();
 sg13g2_fill_2 FILLER_42_24 ();
 sg13g2_decap_8 FILLER_42_48 ();
 sg13g2_decap_4 FILLER_42_55 ();
 sg13g2_decap_8 FILLER_42_78 ();
 sg13g2_fill_1 FILLER_42_85 ();
 sg13g2_fill_2 FILLER_42_101 ();
 sg13g2_fill_2 FILLER_42_108 ();
 sg13g2_fill_1 FILLER_42_142 ();
 sg13g2_decap_8 FILLER_42_191 ();
 sg13g2_fill_2 FILLER_42_198 ();
 sg13g2_fill_1 FILLER_42_200 ();
 sg13g2_fill_1 FILLER_42_205 ();
 sg13g2_decap_8 FILLER_42_215 ();
 sg13g2_decap_4 FILLER_42_222 ();
 sg13g2_fill_2 FILLER_42_226 ();
 sg13g2_fill_2 FILLER_42_232 ();
 sg13g2_fill_1 FILLER_42_234 ();
 sg13g2_decap_4 FILLER_42_250 ();
 sg13g2_fill_2 FILLER_42_254 ();
 sg13g2_decap_4 FILLER_42_259 ();
 sg13g2_fill_1 FILLER_42_263 ();
 sg13g2_decap_4 FILLER_42_318 ();
 sg13g2_decap_8 FILLER_42_342 ();
 sg13g2_decap_8 FILLER_42_349 ();
 sg13g2_fill_2 FILLER_42_356 ();
 sg13g2_fill_2 FILLER_42_401 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_fill_1 FILLER_42_414 ();
 sg13g2_fill_1 FILLER_42_431 ();
 sg13g2_fill_1 FILLER_42_458 ();
 sg13g2_decap_8 FILLER_42_474 ();
 sg13g2_fill_2 FILLER_42_481 ();
 sg13g2_decap_4 FILLER_42_498 ();
 sg13g2_fill_2 FILLER_42_502 ();
 sg13g2_fill_2 FILLER_42_509 ();
 sg13g2_decap_8 FILLER_42_524 ();
 sg13g2_fill_1 FILLER_42_531 ();
 sg13g2_decap_8 FILLER_42_536 ();
 sg13g2_fill_2 FILLER_42_555 ();
 sg13g2_decap_8 FILLER_42_562 ();
 sg13g2_decap_4 FILLER_42_569 ();
 sg13g2_fill_1 FILLER_42_573 ();
 sg13g2_fill_1 FILLER_42_597 ();
 sg13g2_fill_2 FILLER_42_626 ();
 sg13g2_fill_1 FILLER_42_628 ();
 sg13g2_fill_1 FILLER_42_657 ();
 sg13g2_decap_4 FILLER_42_693 ();
 sg13g2_fill_1 FILLER_42_702 ();
 sg13g2_decap_4 FILLER_42_743 ();
 sg13g2_fill_2 FILLER_42_770 ();
 sg13g2_fill_1 FILLER_42_772 ();
 sg13g2_fill_2 FILLER_42_778 ();
 sg13g2_decap_8 FILLER_42_783 ();
 sg13g2_fill_2 FILLER_42_790 ();
 sg13g2_fill_1 FILLER_42_792 ();
 sg13g2_fill_1 FILLER_42_812 ();
 sg13g2_fill_2 FILLER_42_825 ();
 sg13g2_decap_8 FILLER_42_859 ();
 sg13g2_decap_8 FILLER_42_866 ();
 sg13g2_decap_8 FILLER_42_873 ();
 sg13g2_decap_8 FILLER_42_880 ();
 sg13g2_decap_8 FILLER_42_887 ();
 sg13g2_decap_8 FILLER_42_894 ();
 sg13g2_decap_8 FILLER_42_901 ();
 sg13g2_decap_8 FILLER_42_908 ();
 sg13g2_decap_8 FILLER_42_915 ();
 sg13g2_decap_8 FILLER_42_922 ();
 sg13g2_decap_8 FILLER_42_929 ();
 sg13g2_decap_8 FILLER_42_936 ();
 sg13g2_decap_8 FILLER_42_943 ();
 sg13g2_decap_8 FILLER_42_950 ();
 sg13g2_decap_8 FILLER_42_957 ();
 sg13g2_decap_8 FILLER_42_964 ();
 sg13g2_decap_8 FILLER_42_971 ();
 sg13g2_decap_8 FILLER_42_978 ();
 sg13g2_decap_8 FILLER_42_985 ();
 sg13g2_decap_8 FILLER_42_992 ();
 sg13g2_decap_8 FILLER_42_999 ();
 sg13g2_decap_8 FILLER_42_1006 ();
 sg13g2_decap_8 FILLER_42_1013 ();
 sg13g2_decap_8 FILLER_42_1020 ();
 sg13g2_fill_2 FILLER_42_1027 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_decap_4 FILLER_43_55 ();
 sg13g2_fill_2 FILLER_43_59 ();
 sg13g2_decap_8 FILLER_43_76 ();
 sg13g2_decap_8 FILLER_43_83 ();
 sg13g2_decap_4 FILLER_43_90 ();
 sg13g2_fill_1 FILLER_43_94 ();
 sg13g2_decap_8 FILLER_43_107 ();
 sg13g2_decap_4 FILLER_43_130 ();
 sg13g2_decap_4 FILLER_43_143 ();
 sg13g2_fill_1 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_153 ();
 sg13g2_decap_8 FILLER_43_178 ();
 sg13g2_fill_1 FILLER_43_185 ();
 sg13g2_fill_2 FILLER_43_223 ();
 sg13g2_fill_1 FILLER_43_225 ();
 sg13g2_fill_1 FILLER_43_261 ();
 sg13g2_fill_2 FILLER_43_267 ();
 sg13g2_fill_1 FILLER_43_269 ();
 sg13g2_decap_4 FILLER_43_277 ();
 sg13g2_fill_2 FILLER_43_281 ();
 sg13g2_decap_4 FILLER_43_292 ();
 sg13g2_fill_1 FILLER_43_296 ();
 sg13g2_decap_8 FILLER_43_314 ();
 sg13g2_fill_2 FILLER_43_321 ();
 sg13g2_fill_1 FILLER_43_343 ();
 sg13g2_decap_4 FILLER_43_357 ();
 sg13g2_decap_4 FILLER_43_374 ();
 sg13g2_fill_2 FILLER_43_383 ();
 sg13g2_fill_1 FILLER_43_385 ();
 sg13g2_decap_4 FILLER_43_391 ();
 sg13g2_fill_1 FILLER_43_395 ();
 sg13g2_decap_8 FILLER_43_400 ();
 sg13g2_decap_8 FILLER_43_448 ();
 sg13g2_decap_4 FILLER_43_455 ();
 sg13g2_fill_1 FILLER_43_459 ();
 sg13g2_decap_8 FILLER_43_478 ();
 sg13g2_decap_8 FILLER_43_485 ();
 sg13g2_fill_2 FILLER_43_492 ();
 sg13g2_decap_8 FILLER_43_525 ();
 sg13g2_decap_4 FILLER_43_532 ();
 sg13g2_fill_2 FILLER_43_565 ();
 sg13g2_fill_2 FILLER_43_589 ();
 sg13g2_fill_1 FILLER_43_591 ();
 sg13g2_decap_4 FILLER_43_604 ();
 sg13g2_decap_8 FILLER_43_621 ();
 sg13g2_decap_4 FILLER_43_628 ();
 sg13g2_fill_1 FILLER_43_632 ();
 sg13g2_decap_8 FILLER_43_653 ();
 sg13g2_decap_8 FILLER_43_660 ();
 sg13g2_fill_2 FILLER_43_677 ();
 sg13g2_decap_8 FILLER_43_688 ();
 sg13g2_decap_4 FILLER_43_695 ();
 sg13g2_fill_2 FILLER_43_718 ();
 sg13g2_decap_8 FILLER_43_737 ();
 sg13g2_fill_1 FILLER_43_784 ();
 sg13g2_decap_8 FILLER_43_818 ();
 sg13g2_decap_4 FILLER_43_825 ();
 sg13g2_decap_8 FILLER_43_842 ();
 sg13g2_decap_8 FILLER_43_849 ();
 sg13g2_decap_8 FILLER_43_856 ();
 sg13g2_decap_8 FILLER_43_863 ();
 sg13g2_decap_8 FILLER_43_870 ();
 sg13g2_decap_8 FILLER_43_877 ();
 sg13g2_decap_8 FILLER_43_884 ();
 sg13g2_decap_8 FILLER_43_891 ();
 sg13g2_decap_8 FILLER_43_898 ();
 sg13g2_decap_8 FILLER_43_905 ();
 sg13g2_decap_8 FILLER_43_912 ();
 sg13g2_decap_8 FILLER_43_919 ();
 sg13g2_decap_8 FILLER_43_926 ();
 sg13g2_decap_8 FILLER_43_933 ();
 sg13g2_decap_8 FILLER_43_940 ();
 sg13g2_decap_8 FILLER_43_947 ();
 sg13g2_decap_8 FILLER_43_954 ();
 sg13g2_decap_8 FILLER_43_961 ();
 sg13g2_decap_8 FILLER_43_968 ();
 sg13g2_decap_8 FILLER_43_975 ();
 sg13g2_decap_8 FILLER_43_982 ();
 sg13g2_decap_8 FILLER_43_989 ();
 sg13g2_decap_8 FILLER_43_996 ();
 sg13g2_decap_8 FILLER_43_1003 ();
 sg13g2_decap_8 FILLER_43_1010 ();
 sg13g2_decap_8 FILLER_43_1017 ();
 sg13g2_decap_4 FILLER_43_1024 ();
 sg13g2_fill_1 FILLER_43_1028 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_7 ();
 sg13g2_fill_1 FILLER_44_35 ();
 sg13g2_fill_1 FILLER_44_76 ();
 sg13g2_decap_4 FILLER_44_87 ();
 sg13g2_decap_8 FILLER_44_118 ();
 sg13g2_fill_2 FILLER_44_125 ();
 sg13g2_fill_1 FILLER_44_127 ();
 sg13g2_fill_2 FILLER_44_141 ();
 sg13g2_fill_2 FILLER_44_166 ();
 sg13g2_fill_2 FILLER_44_173 ();
 sg13g2_fill_1 FILLER_44_175 ();
 sg13g2_fill_2 FILLER_44_186 ();
 sg13g2_decap_8 FILLER_44_193 ();
 sg13g2_fill_2 FILLER_44_204 ();
 sg13g2_fill_1 FILLER_44_206 ();
 sg13g2_decap_8 FILLER_44_220 ();
 sg13g2_fill_2 FILLER_44_227 ();
 sg13g2_fill_2 FILLER_44_236 ();
 sg13g2_fill_1 FILLER_44_238 ();
 sg13g2_decap_8 FILLER_44_249 ();
 sg13g2_decap_8 FILLER_44_256 ();
 sg13g2_fill_2 FILLER_44_263 ();
 sg13g2_decap_8 FILLER_44_270 ();
 sg13g2_decap_8 FILLER_44_277 ();
 sg13g2_fill_2 FILLER_44_284 ();
 sg13g2_fill_2 FILLER_44_311 ();
 sg13g2_fill_1 FILLER_44_313 ();
 sg13g2_decap_4 FILLER_44_319 ();
 sg13g2_fill_2 FILLER_44_323 ();
 sg13g2_fill_2 FILLER_44_330 ();
 sg13g2_decap_8 FILLER_44_341 ();
 sg13g2_decap_8 FILLER_44_348 ();
 sg13g2_fill_1 FILLER_44_355 ();
 sg13g2_decap_8 FILLER_44_426 ();
 sg13g2_decap_8 FILLER_44_442 ();
 sg13g2_decap_4 FILLER_44_449 ();
 sg13g2_fill_2 FILLER_44_453 ();
 sg13g2_decap_4 FILLER_44_481 ();
 sg13g2_fill_2 FILLER_44_485 ();
 sg13g2_fill_2 FILLER_44_517 ();
 sg13g2_fill_1 FILLER_44_519 ();
 sg13g2_decap_8 FILLER_44_529 ();
 sg13g2_decap_4 FILLER_44_536 ();
 sg13g2_fill_2 FILLER_44_540 ();
 sg13g2_fill_1 FILLER_44_547 ();
 sg13g2_fill_2 FILLER_44_587 ();
 sg13g2_decap_8 FILLER_44_631 ();
 sg13g2_fill_2 FILLER_44_638 ();
 sg13g2_fill_1 FILLER_44_640 ();
 sg13g2_fill_1 FILLER_44_649 ();
 sg13g2_decap_8 FILLER_44_655 ();
 sg13g2_decap_4 FILLER_44_671 ();
 sg13g2_fill_2 FILLER_44_675 ();
 sg13g2_decap_8 FILLER_44_708 ();
 sg13g2_decap_8 FILLER_44_715 ();
 sg13g2_fill_2 FILLER_44_722 ();
 sg13g2_fill_1 FILLER_44_724 ();
 sg13g2_decap_8 FILLER_44_752 ();
 sg13g2_fill_1 FILLER_44_759 ();
 sg13g2_decap_4 FILLER_44_769 ();
 sg13g2_fill_2 FILLER_44_773 ();
 sg13g2_decap_4 FILLER_44_784 ();
 sg13g2_fill_2 FILLER_44_788 ();
 sg13g2_decap_8 FILLER_44_794 ();
 sg13g2_decap_8 FILLER_44_801 ();
 sg13g2_decap_8 FILLER_44_808 ();
 sg13g2_decap_8 FILLER_44_815 ();
 sg13g2_decap_8 FILLER_44_822 ();
 sg13g2_decap_8 FILLER_44_829 ();
 sg13g2_decap_8 FILLER_44_836 ();
 sg13g2_decap_8 FILLER_44_843 ();
 sg13g2_decap_8 FILLER_44_850 ();
 sg13g2_decap_8 FILLER_44_857 ();
 sg13g2_decap_8 FILLER_44_864 ();
 sg13g2_decap_8 FILLER_44_871 ();
 sg13g2_decap_8 FILLER_44_878 ();
 sg13g2_decap_8 FILLER_44_885 ();
 sg13g2_decap_8 FILLER_44_892 ();
 sg13g2_decap_8 FILLER_44_899 ();
 sg13g2_decap_8 FILLER_44_906 ();
 sg13g2_decap_8 FILLER_44_913 ();
 sg13g2_decap_8 FILLER_44_920 ();
 sg13g2_decap_8 FILLER_44_927 ();
 sg13g2_decap_8 FILLER_44_934 ();
 sg13g2_decap_8 FILLER_44_941 ();
 sg13g2_decap_8 FILLER_44_948 ();
 sg13g2_decap_8 FILLER_44_955 ();
 sg13g2_decap_8 FILLER_44_962 ();
 sg13g2_decap_8 FILLER_44_969 ();
 sg13g2_decap_8 FILLER_44_976 ();
 sg13g2_decap_8 FILLER_44_983 ();
 sg13g2_decap_8 FILLER_44_990 ();
 sg13g2_decap_8 FILLER_44_997 ();
 sg13g2_decap_8 FILLER_44_1004 ();
 sg13g2_decap_8 FILLER_44_1011 ();
 sg13g2_decap_8 FILLER_44_1018 ();
 sg13g2_decap_4 FILLER_44_1025 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_12 ();
 sg13g2_decap_4 FILLER_45_17 ();
 sg13g2_fill_2 FILLER_45_30 ();
 sg13g2_fill_1 FILLER_45_32 ();
 sg13g2_decap_8 FILLER_45_50 ();
 sg13g2_fill_2 FILLER_45_57 ();
 sg13g2_fill_1 FILLER_45_59 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_fill_2 FILLER_45_91 ();
 sg13g2_fill_1 FILLER_45_93 ();
 sg13g2_fill_2 FILLER_45_112 ();
 sg13g2_fill_1 FILLER_45_124 ();
 sg13g2_fill_1 FILLER_45_138 ();
 sg13g2_fill_2 FILLER_45_166 ();
 sg13g2_fill_1 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_213 ();
 sg13g2_decap_8 FILLER_45_243 ();
 sg13g2_decap_4 FILLER_45_250 ();
 sg13g2_decap_8 FILLER_45_276 ();
 sg13g2_decap_8 FILLER_45_283 ();
 sg13g2_fill_1 FILLER_45_290 ();
 sg13g2_fill_2 FILLER_45_311 ();
 sg13g2_fill_1 FILLER_45_313 ();
 sg13g2_decap_8 FILLER_45_345 ();
 sg13g2_decap_8 FILLER_45_352 ();
 sg13g2_decap_8 FILLER_45_359 ();
 sg13g2_decap_8 FILLER_45_366 ();
 sg13g2_fill_1 FILLER_45_373 ();
 sg13g2_fill_1 FILLER_45_396 ();
 sg13g2_fill_2 FILLER_45_420 ();
 sg13g2_fill_1 FILLER_45_422 ();
 sg13g2_decap_4 FILLER_45_426 ();
 sg13g2_fill_1 FILLER_45_458 ();
 sg13g2_decap_8 FILLER_45_474 ();
 sg13g2_fill_2 FILLER_45_481 ();
 sg13g2_fill_1 FILLER_45_483 ();
 sg13g2_fill_2 FILLER_45_542 ();
 sg13g2_fill_1 FILLER_45_544 ();
 sg13g2_decap_8 FILLER_45_550 ();
 sg13g2_fill_1 FILLER_45_557 ();
 sg13g2_fill_2 FILLER_45_567 ();
 sg13g2_fill_2 FILLER_45_583 ();
 sg13g2_fill_1 FILLER_45_585 ();
 sg13g2_fill_1 FILLER_45_614 ();
 sg13g2_decap_8 FILLER_45_675 ();
 sg13g2_decap_4 FILLER_45_682 ();
 sg13g2_decap_8 FILLER_45_690 ();
 sg13g2_decap_8 FILLER_45_697 ();
 sg13g2_decap_8 FILLER_45_704 ();
 sg13g2_decap_8 FILLER_45_711 ();
 sg13g2_decap_8 FILLER_45_718 ();
 sg13g2_decap_8 FILLER_45_725 ();
 sg13g2_decap_8 FILLER_45_732 ();
 sg13g2_decap_8 FILLER_45_739 ();
 sg13g2_decap_8 FILLER_45_746 ();
 sg13g2_decap_8 FILLER_45_753 ();
 sg13g2_decap_8 FILLER_45_760 ();
 sg13g2_decap_8 FILLER_45_767 ();
 sg13g2_decap_8 FILLER_45_774 ();
 sg13g2_decap_8 FILLER_45_781 ();
 sg13g2_decap_8 FILLER_45_788 ();
 sg13g2_decap_8 FILLER_45_795 ();
 sg13g2_decap_8 FILLER_45_802 ();
 sg13g2_decap_8 FILLER_45_809 ();
 sg13g2_decap_8 FILLER_45_816 ();
 sg13g2_decap_8 FILLER_45_823 ();
 sg13g2_decap_8 FILLER_45_830 ();
 sg13g2_decap_8 FILLER_45_837 ();
 sg13g2_decap_8 FILLER_45_844 ();
 sg13g2_decap_8 FILLER_45_851 ();
 sg13g2_decap_8 FILLER_45_858 ();
 sg13g2_decap_8 FILLER_45_865 ();
 sg13g2_decap_8 FILLER_45_872 ();
 sg13g2_decap_8 FILLER_45_879 ();
 sg13g2_decap_8 FILLER_45_886 ();
 sg13g2_decap_8 FILLER_45_893 ();
 sg13g2_decap_8 FILLER_45_900 ();
 sg13g2_decap_8 FILLER_45_907 ();
 sg13g2_decap_8 FILLER_45_914 ();
 sg13g2_decap_8 FILLER_45_921 ();
 sg13g2_decap_8 FILLER_45_928 ();
 sg13g2_decap_8 FILLER_45_935 ();
 sg13g2_decap_8 FILLER_45_942 ();
 sg13g2_decap_8 FILLER_45_949 ();
 sg13g2_decap_8 FILLER_45_956 ();
 sg13g2_decap_8 FILLER_45_963 ();
 sg13g2_decap_8 FILLER_45_970 ();
 sg13g2_decap_8 FILLER_45_977 ();
 sg13g2_decap_8 FILLER_45_984 ();
 sg13g2_decap_8 FILLER_45_991 ();
 sg13g2_decap_8 FILLER_45_998 ();
 sg13g2_decap_8 FILLER_45_1005 ();
 sg13g2_decap_8 FILLER_45_1012 ();
 sg13g2_decap_8 FILLER_45_1019 ();
 sg13g2_fill_2 FILLER_45_1026 ();
 sg13g2_fill_1 FILLER_45_1028 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_2 ();
 sg13g2_decap_8 FILLER_46_44 ();
 sg13g2_decap_8 FILLER_46_51 ();
 sg13g2_fill_2 FILLER_46_83 ();
 sg13g2_decap_8 FILLER_46_94 ();
 sg13g2_decap_4 FILLER_46_101 ();
 sg13g2_fill_2 FILLER_46_105 ();
 sg13g2_decap_4 FILLER_46_144 ();
 sg13g2_fill_1 FILLER_46_148 ();
 sg13g2_decap_4 FILLER_46_175 ();
 sg13g2_fill_2 FILLER_46_203 ();
 sg13g2_decap_4 FILLER_46_214 ();
 sg13g2_fill_2 FILLER_46_218 ();
 sg13g2_fill_2 FILLER_46_249 ();
 sg13g2_fill_1 FILLER_46_251 ();
 sg13g2_fill_2 FILLER_46_280 ();
 sg13g2_fill_1 FILLER_46_295 ();
 sg13g2_fill_1 FILLER_46_353 ();
 sg13g2_decap_8 FILLER_46_367 ();
 sg13g2_decap_4 FILLER_46_374 ();
 sg13g2_fill_1 FILLER_46_378 ();
 sg13g2_decap_8 FILLER_46_398 ();
 sg13g2_decap_8 FILLER_46_405 ();
 sg13g2_fill_2 FILLER_46_412 ();
 sg13g2_fill_1 FILLER_46_414 ();
 sg13g2_decap_4 FILLER_46_418 ();
 sg13g2_decap_8 FILLER_46_450 ();
 sg13g2_decap_4 FILLER_46_457 ();
 sg13g2_fill_2 FILLER_46_461 ();
 sg13g2_decap_4 FILLER_46_470 ();
 sg13g2_fill_2 FILLER_46_483 ();
 sg13g2_fill_1 FILLER_46_485 ();
 sg13g2_fill_1 FILLER_46_494 ();
 sg13g2_decap_8 FILLER_46_527 ();
 sg13g2_decap_8 FILLER_46_534 ();
 sg13g2_decap_8 FILLER_46_546 ();
 sg13g2_decap_4 FILLER_46_553 ();
 sg13g2_fill_1 FILLER_46_557 ();
 sg13g2_decap_8 FILLER_46_620 ();
 sg13g2_fill_1 FILLER_46_631 ();
 sg13g2_decap_8 FILLER_46_641 ();
 sg13g2_decap_4 FILLER_46_648 ();
 sg13g2_decap_8 FILLER_46_656 ();
 sg13g2_decap_8 FILLER_46_663 ();
 sg13g2_decap_8 FILLER_46_670 ();
 sg13g2_decap_8 FILLER_46_677 ();
 sg13g2_decap_8 FILLER_46_684 ();
 sg13g2_decap_8 FILLER_46_691 ();
 sg13g2_decap_8 FILLER_46_698 ();
 sg13g2_decap_8 FILLER_46_705 ();
 sg13g2_decap_8 FILLER_46_712 ();
 sg13g2_decap_8 FILLER_46_719 ();
 sg13g2_decap_8 FILLER_46_726 ();
 sg13g2_decap_8 FILLER_46_733 ();
 sg13g2_decap_8 FILLER_46_740 ();
 sg13g2_decap_8 FILLER_46_747 ();
 sg13g2_decap_8 FILLER_46_754 ();
 sg13g2_decap_8 FILLER_46_761 ();
 sg13g2_decap_8 FILLER_46_768 ();
 sg13g2_decap_8 FILLER_46_775 ();
 sg13g2_decap_8 FILLER_46_782 ();
 sg13g2_decap_8 FILLER_46_789 ();
 sg13g2_decap_8 FILLER_46_796 ();
 sg13g2_decap_8 FILLER_46_803 ();
 sg13g2_decap_8 FILLER_46_810 ();
 sg13g2_decap_8 FILLER_46_817 ();
 sg13g2_decap_8 FILLER_46_824 ();
 sg13g2_decap_8 FILLER_46_831 ();
 sg13g2_decap_8 FILLER_46_838 ();
 sg13g2_decap_8 FILLER_46_845 ();
 sg13g2_decap_8 FILLER_46_852 ();
 sg13g2_decap_8 FILLER_46_859 ();
 sg13g2_decap_8 FILLER_46_866 ();
 sg13g2_decap_8 FILLER_46_873 ();
 sg13g2_decap_8 FILLER_46_880 ();
 sg13g2_decap_8 FILLER_46_887 ();
 sg13g2_decap_8 FILLER_46_894 ();
 sg13g2_decap_8 FILLER_46_901 ();
 sg13g2_decap_8 FILLER_46_908 ();
 sg13g2_decap_8 FILLER_46_915 ();
 sg13g2_decap_8 FILLER_46_922 ();
 sg13g2_decap_8 FILLER_46_929 ();
 sg13g2_decap_8 FILLER_46_936 ();
 sg13g2_decap_8 FILLER_46_943 ();
 sg13g2_decap_8 FILLER_46_950 ();
 sg13g2_decap_8 FILLER_46_957 ();
 sg13g2_decap_8 FILLER_46_964 ();
 sg13g2_decap_8 FILLER_46_971 ();
 sg13g2_decap_8 FILLER_46_978 ();
 sg13g2_decap_8 FILLER_46_985 ();
 sg13g2_decap_8 FILLER_46_992 ();
 sg13g2_decap_8 FILLER_46_999 ();
 sg13g2_decap_8 FILLER_46_1006 ();
 sg13g2_decap_8 FILLER_46_1013 ();
 sg13g2_decap_8 FILLER_46_1020 ();
 sg13g2_fill_2 FILLER_46_1027 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_fill_2 FILLER_47_28 ();
 sg13g2_fill_1 FILLER_47_30 ();
 sg13g2_fill_1 FILLER_47_62 ();
 sg13g2_fill_1 FILLER_47_96 ();
 sg13g2_fill_1 FILLER_47_111 ();
 sg13g2_fill_2 FILLER_47_120 ();
 sg13g2_decap_4 FILLER_47_149 ();
 sg13g2_fill_1 FILLER_47_153 ();
 sg13g2_fill_1 FILLER_47_164 ();
 sg13g2_fill_1 FILLER_47_179 ();
 sg13g2_fill_2 FILLER_47_189 ();
 sg13g2_fill_2 FILLER_47_222 ();
 sg13g2_decap_4 FILLER_47_251 ();
 sg13g2_fill_2 FILLER_47_255 ();
 sg13g2_fill_2 FILLER_47_280 ();
 sg13g2_decap_4 FILLER_47_317 ();
 sg13g2_decap_4 FILLER_47_330 ();
 sg13g2_fill_1 FILLER_47_334 ();
 sg13g2_decap_8 FILLER_47_340 ();
 sg13g2_fill_2 FILLER_47_347 ();
 sg13g2_fill_2 FILLER_47_377 ();
 sg13g2_fill_1 FILLER_47_379 ();
 sg13g2_decap_8 FILLER_47_407 ();
 sg13g2_decap_8 FILLER_47_414 ();
 sg13g2_decap_4 FILLER_47_421 ();
 sg13g2_decap_8 FILLER_47_442 ();
 sg13g2_decap_8 FILLER_47_449 ();
 sg13g2_decap_4 FILLER_47_456 ();
 sg13g2_fill_1 FILLER_47_460 ();
 sg13g2_decap_8 FILLER_47_489 ();
 sg13g2_decap_4 FILLER_47_496 ();
 sg13g2_decap_8 FILLER_47_504 ();
 sg13g2_decap_8 FILLER_47_520 ();
 sg13g2_decap_8 FILLER_47_527 ();
 sg13g2_decap_4 FILLER_47_534 ();
 sg13g2_fill_2 FILLER_47_565 ();
 sg13g2_decap_8 FILLER_47_571 ();
 sg13g2_decap_8 FILLER_47_578 ();
 sg13g2_decap_4 FILLER_47_585 ();
 sg13g2_fill_2 FILLER_47_589 ();
 sg13g2_decap_8 FILLER_47_595 ();
 sg13g2_decap_4 FILLER_47_602 ();
 sg13g2_fill_2 FILLER_47_606 ();
 sg13g2_decap_8 FILLER_47_612 ();
 sg13g2_decap_8 FILLER_47_619 ();
 sg13g2_decap_8 FILLER_47_626 ();
 sg13g2_decap_8 FILLER_47_633 ();
 sg13g2_decap_8 FILLER_47_640 ();
 sg13g2_decap_8 FILLER_47_647 ();
 sg13g2_decap_8 FILLER_47_654 ();
 sg13g2_decap_8 FILLER_47_661 ();
 sg13g2_decap_8 FILLER_47_668 ();
 sg13g2_decap_8 FILLER_47_675 ();
 sg13g2_decap_8 FILLER_47_682 ();
 sg13g2_decap_8 FILLER_47_689 ();
 sg13g2_decap_8 FILLER_47_696 ();
 sg13g2_decap_8 FILLER_47_703 ();
 sg13g2_decap_8 FILLER_47_710 ();
 sg13g2_decap_8 FILLER_47_717 ();
 sg13g2_decap_8 FILLER_47_724 ();
 sg13g2_decap_8 FILLER_47_731 ();
 sg13g2_decap_8 FILLER_47_738 ();
 sg13g2_decap_8 FILLER_47_745 ();
 sg13g2_decap_8 FILLER_47_752 ();
 sg13g2_decap_8 FILLER_47_759 ();
 sg13g2_decap_8 FILLER_47_766 ();
 sg13g2_decap_8 FILLER_47_773 ();
 sg13g2_decap_8 FILLER_47_780 ();
 sg13g2_decap_8 FILLER_47_787 ();
 sg13g2_decap_8 FILLER_47_794 ();
 sg13g2_decap_8 FILLER_47_801 ();
 sg13g2_decap_8 FILLER_47_808 ();
 sg13g2_decap_8 FILLER_47_815 ();
 sg13g2_decap_8 FILLER_47_822 ();
 sg13g2_decap_8 FILLER_47_829 ();
 sg13g2_decap_8 FILLER_47_836 ();
 sg13g2_decap_8 FILLER_47_843 ();
 sg13g2_decap_8 FILLER_47_850 ();
 sg13g2_decap_8 FILLER_47_857 ();
 sg13g2_decap_8 FILLER_47_864 ();
 sg13g2_decap_8 FILLER_47_871 ();
 sg13g2_decap_8 FILLER_47_878 ();
 sg13g2_decap_8 FILLER_47_885 ();
 sg13g2_decap_8 FILLER_47_892 ();
 sg13g2_decap_8 FILLER_47_899 ();
 sg13g2_decap_8 FILLER_47_906 ();
 sg13g2_decap_8 FILLER_47_913 ();
 sg13g2_decap_8 FILLER_47_920 ();
 sg13g2_decap_8 FILLER_47_927 ();
 sg13g2_decap_8 FILLER_47_934 ();
 sg13g2_decap_8 FILLER_47_941 ();
 sg13g2_decap_8 FILLER_47_948 ();
 sg13g2_decap_8 FILLER_47_955 ();
 sg13g2_decap_8 FILLER_47_962 ();
 sg13g2_decap_8 FILLER_47_969 ();
 sg13g2_decap_8 FILLER_47_976 ();
 sg13g2_decap_8 FILLER_47_983 ();
 sg13g2_decap_8 FILLER_47_990 ();
 sg13g2_decap_8 FILLER_47_997 ();
 sg13g2_decap_8 FILLER_47_1004 ();
 sg13g2_decap_8 FILLER_47_1011 ();
 sg13g2_decap_8 FILLER_47_1018 ();
 sg13g2_decap_4 FILLER_47_1025 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_4 FILLER_48_35 ();
 sg13g2_fill_1 FILLER_48_39 ();
 sg13g2_fill_2 FILLER_48_44 ();
 sg13g2_fill_1 FILLER_48_46 ();
 sg13g2_fill_2 FILLER_48_130 ();
 sg13g2_fill_1 FILLER_48_132 ();
 sg13g2_decap_4 FILLER_48_205 ();
 sg13g2_fill_1 FILLER_48_209 ();
 sg13g2_decap_4 FILLER_48_294 ();
 sg13g2_fill_2 FILLER_48_363 ();
 sg13g2_decap_4 FILLER_48_378 ();
 sg13g2_fill_2 FILLER_48_382 ();
 sg13g2_decap_4 FILLER_48_393 ();
 sg13g2_fill_2 FILLER_48_397 ();
 sg13g2_decap_8 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_48_415 ();
 sg13g2_decap_8 FILLER_48_422 ();
 sg13g2_decap_8 FILLER_48_429 ();
 sg13g2_decap_8 FILLER_48_436 ();
 sg13g2_decap_8 FILLER_48_443 ();
 sg13g2_decap_8 FILLER_48_450 ();
 sg13g2_decap_8 FILLER_48_457 ();
 sg13g2_decap_8 FILLER_48_464 ();
 sg13g2_decap_8 FILLER_48_471 ();
 sg13g2_decap_8 FILLER_48_478 ();
 sg13g2_decap_8 FILLER_48_485 ();
 sg13g2_decap_8 FILLER_48_492 ();
 sg13g2_decap_8 FILLER_48_499 ();
 sg13g2_decap_8 FILLER_48_506 ();
 sg13g2_decap_8 FILLER_48_513 ();
 sg13g2_decap_8 FILLER_48_520 ();
 sg13g2_decap_8 FILLER_48_527 ();
 sg13g2_decap_8 FILLER_48_534 ();
 sg13g2_fill_2 FILLER_48_541 ();
 sg13g2_decap_8 FILLER_48_547 ();
 sg13g2_decap_8 FILLER_48_563 ();
 sg13g2_decap_8 FILLER_48_570 ();
 sg13g2_decap_8 FILLER_48_577 ();
 sg13g2_decap_8 FILLER_48_584 ();
 sg13g2_decap_8 FILLER_48_591 ();
 sg13g2_decap_8 FILLER_48_598 ();
 sg13g2_decap_8 FILLER_48_605 ();
 sg13g2_decap_8 FILLER_48_612 ();
 sg13g2_decap_8 FILLER_48_619 ();
 sg13g2_decap_8 FILLER_48_626 ();
 sg13g2_decap_8 FILLER_48_633 ();
 sg13g2_decap_8 FILLER_48_640 ();
 sg13g2_decap_8 FILLER_48_647 ();
 sg13g2_decap_8 FILLER_48_654 ();
 sg13g2_decap_8 FILLER_48_661 ();
 sg13g2_decap_8 FILLER_48_668 ();
 sg13g2_decap_8 FILLER_48_675 ();
 sg13g2_decap_8 FILLER_48_682 ();
 sg13g2_decap_8 FILLER_48_689 ();
 sg13g2_decap_8 FILLER_48_696 ();
 sg13g2_decap_8 FILLER_48_703 ();
 sg13g2_decap_8 FILLER_48_710 ();
 sg13g2_decap_8 FILLER_48_717 ();
 sg13g2_decap_8 FILLER_48_724 ();
 sg13g2_decap_8 FILLER_48_731 ();
 sg13g2_decap_8 FILLER_48_738 ();
 sg13g2_decap_8 FILLER_48_745 ();
 sg13g2_decap_8 FILLER_48_752 ();
 sg13g2_decap_8 FILLER_48_759 ();
 sg13g2_decap_8 FILLER_48_766 ();
 sg13g2_decap_8 FILLER_48_773 ();
 sg13g2_decap_8 FILLER_48_780 ();
 sg13g2_decap_8 FILLER_48_787 ();
 sg13g2_decap_8 FILLER_48_794 ();
 sg13g2_decap_8 FILLER_48_801 ();
 sg13g2_decap_8 FILLER_48_808 ();
 sg13g2_decap_8 FILLER_48_815 ();
 sg13g2_decap_8 FILLER_48_822 ();
 sg13g2_decap_8 FILLER_48_829 ();
 sg13g2_decap_8 FILLER_48_836 ();
 sg13g2_decap_8 FILLER_48_843 ();
 sg13g2_decap_8 FILLER_48_850 ();
 sg13g2_decap_8 FILLER_48_857 ();
 sg13g2_decap_8 FILLER_48_864 ();
 sg13g2_decap_8 FILLER_48_871 ();
 sg13g2_decap_8 FILLER_48_878 ();
 sg13g2_decap_8 FILLER_48_885 ();
 sg13g2_decap_8 FILLER_48_892 ();
 sg13g2_decap_8 FILLER_48_899 ();
 sg13g2_decap_8 FILLER_48_906 ();
 sg13g2_decap_8 FILLER_48_913 ();
 sg13g2_decap_8 FILLER_48_920 ();
 sg13g2_decap_8 FILLER_48_927 ();
 sg13g2_decap_8 FILLER_48_934 ();
 sg13g2_decap_8 FILLER_48_941 ();
 sg13g2_decap_8 FILLER_48_948 ();
 sg13g2_decap_8 FILLER_48_955 ();
 sg13g2_decap_8 FILLER_48_962 ();
 sg13g2_decap_8 FILLER_48_969 ();
 sg13g2_decap_8 FILLER_48_976 ();
 sg13g2_decap_8 FILLER_48_983 ();
 sg13g2_decap_8 FILLER_48_990 ();
 sg13g2_decap_8 FILLER_48_997 ();
 sg13g2_decap_8 FILLER_48_1004 ();
 sg13g2_decap_8 FILLER_48_1011 ();
 sg13g2_decap_8 FILLER_48_1018 ();
 sg13g2_decap_4 FILLER_48_1025 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_fill_2 FILLER_49_49 ();
 sg13g2_fill_1 FILLER_49_51 ();
 sg13g2_fill_2 FILLER_49_59 ();
 sg13g2_fill_1 FILLER_49_61 ();
 sg13g2_fill_2 FILLER_49_80 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_4 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_134 ();
 sg13g2_fill_2 FILLER_49_141 ();
 sg13g2_decap_8 FILLER_49_160 ();
 sg13g2_decap_8 FILLER_49_167 ();
 sg13g2_decap_4 FILLER_49_174 ();
 sg13g2_decap_8 FILLER_49_182 ();
 sg13g2_decap_8 FILLER_49_189 ();
 sg13g2_decap_8 FILLER_49_196 ();
 sg13g2_decap_8 FILLER_49_203 ();
 sg13g2_decap_8 FILLER_49_210 ();
 sg13g2_fill_2 FILLER_49_217 ();
 sg13g2_fill_1 FILLER_49_219 ();
 sg13g2_decap_8 FILLER_49_227 ();
 sg13g2_decap_8 FILLER_49_234 ();
 sg13g2_decap_8 FILLER_49_241 ();
 sg13g2_decap_8 FILLER_49_252 ();
 sg13g2_decap_8 FILLER_49_259 ();
 sg13g2_decap_4 FILLER_49_266 ();
 sg13g2_fill_1 FILLER_49_270 ();
 sg13g2_decap_8 FILLER_49_275 ();
 sg13g2_fill_2 FILLER_49_282 ();
 sg13g2_decap_8 FILLER_49_297 ();
 sg13g2_decap_8 FILLER_49_304 ();
 sg13g2_fill_2 FILLER_49_311 ();
 sg13g2_fill_1 FILLER_49_313 ();
 sg13g2_decap_8 FILLER_49_318 ();
 sg13g2_decap_8 FILLER_49_325 ();
 sg13g2_decap_4 FILLER_49_332 ();
 sg13g2_fill_1 FILLER_49_339 ();
 sg13g2_decap_4 FILLER_49_344 ();
 sg13g2_fill_2 FILLER_49_348 ();
 sg13g2_decap_8 FILLER_49_359 ();
 sg13g2_decap_8 FILLER_49_366 ();
 sg13g2_decap_8 FILLER_49_373 ();
 sg13g2_decap_8 FILLER_49_380 ();
 sg13g2_decap_8 FILLER_49_387 ();
 sg13g2_decap_8 FILLER_49_394 ();
 sg13g2_decap_8 FILLER_49_401 ();
 sg13g2_decap_8 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_49_415 ();
 sg13g2_decap_8 FILLER_49_422 ();
 sg13g2_decap_8 FILLER_49_429 ();
 sg13g2_decap_8 FILLER_49_436 ();
 sg13g2_decap_8 FILLER_49_443 ();
 sg13g2_decap_8 FILLER_49_450 ();
 sg13g2_decap_8 FILLER_49_457 ();
 sg13g2_decap_8 FILLER_49_464 ();
 sg13g2_decap_8 FILLER_49_471 ();
 sg13g2_decap_8 FILLER_49_478 ();
 sg13g2_decap_8 FILLER_49_485 ();
 sg13g2_decap_8 FILLER_49_492 ();
 sg13g2_decap_8 FILLER_49_499 ();
 sg13g2_decap_8 FILLER_49_506 ();
 sg13g2_decap_8 FILLER_49_513 ();
 sg13g2_decap_8 FILLER_49_520 ();
 sg13g2_decap_8 FILLER_49_527 ();
 sg13g2_decap_8 FILLER_49_534 ();
 sg13g2_decap_8 FILLER_49_541 ();
 sg13g2_decap_8 FILLER_49_548 ();
 sg13g2_decap_8 FILLER_49_555 ();
 sg13g2_decap_8 FILLER_49_562 ();
 sg13g2_decap_8 FILLER_49_569 ();
 sg13g2_decap_8 FILLER_49_576 ();
 sg13g2_decap_8 FILLER_49_583 ();
 sg13g2_decap_8 FILLER_49_590 ();
 sg13g2_decap_8 FILLER_49_597 ();
 sg13g2_decap_8 FILLER_49_604 ();
 sg13g2_decap_8 FILLER_49_611 ();
 sg13g2_decap_8 FILLER_49_618 ();
 sg13g2_decap_8 FILLER_49_625 ();
 sg13g2_decap_8 FILLER_49_632 ();
 sg13g2_decap_8 FILLER_49_639 ();
 sg13g2_decap_8 FILLER_49_646 ();
 sg13g2_decap_8 FILLER_49_653 ();
 sg13g2_decap_8 FILLER_49_660 ();
 sg13g2_decap_8 FILLER_49_667 ();
 sg13g2_decap_8 FILLER_49_674 ();
 sg13g2_decap_8 FILLER_49_681 ();
 sg13g2_decap_8 FILLER_49_688 ();
 sg13g2_decap_8 FILLER_49_695 ();
 sg13g2_decap_8 FILLER_49_702 ();
 sg13g2_decap_8 FILLER_49_709 ();
 sg13g2_decap_8 FILLER_49_716 ();
 sg13g2_decap_8 FILLER_49_723 ();
 sg13g2_decap_8 FILLER_49_730 ();
 sg13g2_decap_8 FILLER_49_737 ();
 sg13g2_decap_8 FILLER_49_744 ();
 sg13g2_decap_8 FILLER_49_751 ();
 sg13g2_decap_8 FILLER_49_758 ();
 sg13g2_decap_8 FILLER_49_765 ();
 sg13g2_decap_8 FILLER_49_772 ();
 sg13g2_decap_8 FILLER_49_779 ();
 sg13g2_decap_8 FILLER_49_786 ();
 sg13g2_decap_8 FILLER_49_793 ();
 sg13g2_decap_8 FILLER_49_800 ();
 sg13g2_decap_8 FILLER_49_807 ();
 sg13g2_decap_8 FILLER_49_814 ();
 sg13g2_decap_8 FILLER_49_821 ();
 sg13g2_decap_8 FILLER_49_828 ();
 sg13g2_decap_8 FILLER_49_835 ();
 sg13g2_decap_8 FILLER_49_842 ();
 sg13g2_decap_8 FILLER_49_849 ();
 sg13g2_decap_8 FILLER_49_856 ();
 sg13g2_decap_8 FILLER_49_863 ();
 sg13g2_decap_8 FILLER_49_870 ();
 sg13g2_decap_8 FILLER_49_877 ();
 sg13g2_decap_8 FILLER_49_884 ();
 sg13g2_decap_8 FILLER_49_891 ();
 sg13g2_decap_8 FILLER_49_898 ();
 sg13g2_decap_8 FILLER_49_905 ();
 sg13g2_decap_8 FILLER_49_912 ();
 sg13g2_decap_8 FILLER_49_919 ();
 sg13g2_decap_8 FILLER_49_926 ();
 sg13g2_decap_8 FILLER_49_933 ();
 sg13g2_decap_8 FILLER_49_940 ();
 sg13g2_decap_8 FILLER_49_947 ();
 sg13g2_decap_8 FILLER_49_954 ();
 sg13g2_decap_8 FILLER_49_961 ();
 sg13g2_decap_8 FILLER_49_968 ();
 sg13g2_decap_8 FILLER_49_975 ();
 sg13g2_decap_8 FILLER_49_982 ();
 sg13g2_decap_8 FILLER_49_989 ();
 sg13g2_decap_8 FILLER_49_996 ();
 sg13g2_decap_8 FILLER_49_1003 ();
 sg13g2_decap_8 FILLER_49_1010 ();
 sg13g2_decap_8 FILLER_49_1017 ();
 sg13g2_decap_4 FILLER_49_1024 ();
 sg13g2_fill_1 FILLER_49_1028 ();
 assign uio_oe[0] = net10;
 assign uio_oe[1] = net11;
 assign uio_oe[2] = net295;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net296;
 assign uio_oe[6] = net14;
 assign uio_oe[7] = net15;
 assign uio_out[0] = net16;
 assign uio_out[1] = net17;
 assign uio_out[3] = net18;
 assign uio_out[4] = net19;
 assign uio_out[5] = net20;
 assign uio_out[6] = net21;
 assign uio_out[7] = net22;
endmodule
