* NGSPICE file created from heichips25_top_sorter.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_inv_8 abstract view
.subckt sg13g2_inv_8 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

.subckt heichips25_top_sorter VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
XFILLER_39_233 VPWR VGND sg13g2_fill_2
X_3155_ _1606_ VPWR _1607_ VGND net1327 net419 sg13g2_o21ai_1
XFILLER_36_973 VPWR VGND sg13g2_decap_8
XFILLER_35_494 VPWR VGND sg13g2_decap_8
X_3988_ _2361_ net946 net348 VPWR VGND sg13g2_nand2_1
X_5727_ net1024 net1075 _1361_ VPWR VGND sg13g2_nor2b_1
X_5658_ s0.data_out\[10\]\[0\] s0.data_out\[9\]\[0\] net1041 _1303_ VPWR VGND sg13g2_mux2_1
X_4609_ _0351_ VPWR _0352_ VGND _0347_ _0350_ sg13g2_o21ai_1
X_5589_ net1035 net1074 _1242_ VPWR VGND sg13g2_nor2b_1
XFILLER_2_549 VPWR VGND sg13g2_decap_8
X_6134__141 VPWR VGND net141 sg13g2_tiehi
XFILLER_19_907 VPWR VGND sg13g2_fill_1
XFILLER_46_726 VPWR VGND sg13g2_decap_8
XFILLER_27_995 VPWR VGND sg13g2_decap_8
XFILLER_42_943 VPWR VGND sg13g2_decap_8
XFILLER_41_453 VPWR VGND sg13g2_fill_2
XFILLER_9_104 VPWR VGND sg13g2_fill_1
XFILLER_14_667 VPWR VGND sg13g2_fill_1
XFILLER_14_678 VPWR VGND sg13g2_decap_8
XFILLER_6_877 VPWR VGND sg13g2_decap_8
XFILLER_5_343 VPWR VGND sg13g2_decap_4
XFILLER_1_571 VPWR VGND sg13g2_decap_8
XFILLER_49_520 VPWR VGND sg13g2_decap_8
XFILLER_49_597 VPWR VGND sg13g2_decap_8
XFILLER_18_973 VPWR VGND sg13g2_decap_8
XFILLER_45_781 VPWR VGND sg13g2_decap_8
X_4960_ _0670_ VPWR _0671_ VGND net1320 net445 sg13g2_o21ai_1
X_4891_ _0608_ net1264 _0607_ VPWR VGND sg13g2_nand2_1
X_3911_ _2292_ net928 _2291_ VPWR VGND sg13g2_nand2_1
X_3842_ VGND VPWR net954 net495 _2228_ _2227_ sg13g2_a21oi_1
XFILLER_33_976 VPWR VGND sg13g2_decap_8
XFILLER_20_648 VPWR VGND sg13g2_fill_1
X_3773_ VGND VPWR net1222 net957 _2168_ _2166_ sg13g2_a21oi_1
XFILLER_9_660 VPWR VGND sg13g2_fill_2
X_5512_ net1344 VPWR _1171_ VGND net939 _1170_ sg13g2_o21ai_1
X_5443_ _1091_ _1092_ _1112_ VPWR VGND sg13g2_nor2b_1
X_5374_ VGND VPWR _1046_ net501 net1336 sg13g2_or2_1
X_4325_ net1286 VPWR _2658_ VGND net931 _2657_ sg13g2_o21ai_1
X_6118__158 VPWR VGND net158 sg13g2_tiehi
X_4256_ s0.data_out\[21\]\[6\] s0.data_out\[20\]\[6\] net1200 _2596_ VPWR VGND sg13g2_mux2_1
XFILLER_41_1024 VPWR VGND sg13g2_decap_4
X_4187_ _2530_ _2532_ net1285 _2533_ VPWR VGND sg13g2_nand3_1
X_3207_ VGND VPWR net1001 _1651_ _1652_ _1611_ sg13g2_a21oi_1
X_3138_ net1329 VPWR _1593_ VGND _1588_ _1590_ sg13g2_o21ai_1
XFILLER_43_718 VPWR VGND sg13g2_fill_2
XFILLER_24_965 VPWR VGND sg13g2_decap_8
XFILLER_10_136 VPWR VGND sg13g2_decap_8
XFILLER_12_10 VPWR VGND sg13g2_fill_1
XFILLER_3_803 VPWR VGND sg13g2_decap_8
Xhold170 _0188_ VPWR VGND net466 sg13g2_dlygate4sd3_1
Xhold181 s0.data_out\[13\]\[2\] VPWR VGND net477 sg13g2_dlygate4sd3_1
Xhold192 s0.data_out\[2\]\[2\] VPWR VGND net488 sg13g2_dlygate4sd3_1
XFILLER_46_534 VPWR VGND sg13g2_decap_8
XFILLER_37_62 VPWR VGND sg13g2_decap_8
XFILLER_34_707 VPWR VGND sg13g2_decap_8
XFILLER_37_95 VPWR VGND sg13g2_decap_8
XFILLER_41_250 VPWR VGND sg13g2_fill_1
XFILLER_15_987 VPWR VGND sg13g2_decap_8
XFILLER_18_1015 VPWR VGND sg13g2_decap_8
XFILLER_41_294 VPWR VGND sg13g2_fill_1
XFILLER_10_670 VPWR VGND sg13g2_decap_4
XFILLER_5_140 VPWR VGND sg13g2_decap_8
X_4110_ VPWR _2469_ net1004 VGND sg13g2_inv_1
X_5090_ net1333 VPWR _0789_ VGND net937 _0788_ sg13g2_o21ai_1
X_4041_ _2407_ VPWR _2408_ VGND net940 _2347_ sg13g2_o21ai_1
XFILLER_49_394 VPWR VGND sg13g2_decap_8
XFILLER_37_567 VPWR VGND sg13g2_fill_1
X_5992_ net294 VGND VPWR _0042_ s0.data_out\[18\]\[3\] clknet_leaf_35_clk sg13g2_dfrbpq_2
XFILLER_18_781 VPWR VGND sg13g2_decap_8
X_4943_ _0652_ _0655_ net1318 _0656_ VPWR VGND sg13g2_nand3_1
XFILLER_21_913 VPWR VGND sg13g2_fill_2
X_4874_ s0.data_out\[16\]\[2\] s0.data_out\[15\]\[2\] net1141 _0591_ VPWR VGND sg13g2_mux2_1
X_3825_ net953 s0.data_out\[1\]\[5\] _2213_ VPWR VGND sg13g2_and2_1
X_3756_ _2152_ net963 _2098_ _2153_ VPWR VGND sg13g2_a21o_1
X_5426_ _1095_ net1097 net330 VPWR VGND sg13g2_nand2_1
X_3687_ VPWR _0229_ net510 VGND sg13g2_inv_1
XFILLER_0_817 VPWR VGND sg13g2_decap_8
X_5357_ net1103 VPWR _1031_ VGND _1029_ _1030_ sg13g2_o21ai_1
X_4308_ net1178 net1069 _2643_ VPWR VGND sg13g2_nor2b_1
X_5288_ _0969_ net1111 net588 VPWR VGND sg13g2_nand2_1
X_4239_ _2578_ net1190 _2514_ _2579_ VPWR VGND sg13g2_a21o_1
X_6131__144 VPWR VGND net144 sg13g2_tiehi
XFILLER_16_729 VPWR VGND sg13g2_fill_1
XFILLER_24_773 VPWR VGND sg13g2_decap_4
XFILLER_11_445 VPWR VGND sg13g2_decap_4
XFILLER_12_957 VPWR VGND sg13g2_decap_8
X_5961__56 VPWR VGND net56 sg13g2_tiehi
XFILLER_20_990 VPWR VGND sg13g2_decap_8
XFILLER_47_843 VPWR VGND sg13g2_decap_8
XFILLER_46_353 VPWR VGND sg13g2_fill_1
XFILLER_9_33 VPWR VGND sg13g2_fill_1
X_4590_ net1158 net1058 _0335_ VPWR VGND sg13g2_nor2b_1
X_3610_ _2018_ VPWR _2019_ VGND _2011_ _2012_ sg13g2_o21ai_1
XFILLER_7_950 VPWR VGND sg13g2_decap_8
X_6078__201 VPWR VGND net201 sg13g2_tiehi
X_3541_ _1956_ VPWR _1957_ VGND net1312 net433 sg13g2_o21ai_1
XFILLER_6_471 VPWR VGND sg13g2_decap_8
X_3472_ VGND VPWR net981 _1892_ _1893_ _1830_ sg13g2_a21oi_1
X_5211_ net1116 VPWR _0899_ VGND _0897_ _0898_ sg13g2_o21ai_1
XFILLER_9_1013 VPWR VGND sg13g2_decap_8
X_6191_ net79 VGND VPWR _0241_ s0.data_out\[2\]\[3\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_5142_ VGND VPWR net1113 _0834_ _0835_ _0774_ sg13g2_a21oi_1
XFILLER_29_0 VPWR VGND sg13g2_fill_2
XFILLER_38_832 VPWR VGND sg13g2_decap_4
X_5073_ net1113 net1075 _0774_ VPWR VGND sg13g2_nor2b_1
X_4024_ net297 net1208 _2396_ _0258_ VPWR VGND sg13g2_nor3_1
XFILLER_37_364 VPWR VGND sg13g2_fill_2
X_5975_ net41 VGND VPWR net324 s0.was_valid_out\[19\][0] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_4926_ net1139 VPWR _0641_ VGND net1228 net1125 sg13g2_o21ai_1
XFILLER_33_570 VPWR VGND sg13g2_fill_2
XFILLER_20_242 VPWR VGND sg13g2_decap_8
X_4857_ VPWR _0068_ _0576_ VGND sg13g2_inv_1
X_3808_ _2198_ net930 _2197_ VPWR VGND sg13g2_nand2_1
XFILLER_5_909 VPWR VGND sg13g2_decap_8
X_4788_ _0517_ net1214 _0511_ VPWR VGND sg13g2_xnor2_1
X_3739_ _2136_ net966 net553 VPWR VGND sg13g2_nand2_1
X_5409_ _1077_ VPWR _1078_ VGND net1096 _2488_ sg13g2_o21ai_1
XFILLER_0_614 VPWR VGND sg13g2_decap_8
XFILLER_29_843 VPWR VGND sg13g2_fill_2
XFILLER_44_857 VPWR VGND sg13g2_decap_8
XFILLER_34_41 VPWR VGND sg13g2_fill_2
XFILLER_12_754 VPWR VGND sg13g2_fill_2
XFILLER_4_942 VPWR VGND sg13g2_decap_8
XFILLER_3_485 VPWR VGND sg13g2_decap_8
Xfanout1231 net1234 net1231 VPWR VGND sg13g2_buf_8
Xfanout1220 _2450_ net1220 VPWR VGND sg13g2_buf_8
Xfanout1242 net1245 net1242 VPWR VGND sg13g2_buf_8
Xfanout1253 ui_in[5] net1253 VPWR VGND sg13g2_buf_8
Xfanout1264 net1267 net1264 VPWR VGND sg13g2_buf_8
XFILLER_47_640 VPWR VGND sg13g2_decap_8
Xfanout1286 net1288 net1286 VPWR VGND sg13g2_buf_8
Xfanout1275 net1276 net1275 VPWR VGND sg13g2_buf_8
Xfanout1297 net1300 net1297 VPWR VGND sg13g2_buf_8
XFILLER_34_334 VPWR VGND sg13g2_fill_2
XFILLER_22_507 VPWR VGND sg13g2_decap_8
X_5760_ net1037 VPWR _1390_ VGND _1388_ _1389_ sg13g2_o21ai_1
X_4711_ net1147 net1062 _0445_ VPWR VGND sg13g2_nor2b_1
X_5691_ _1336_ _1331_ _1335_ VPWR VGND sg13g2_nand2_1
X_4642_ _0382_ net1157 _0355_ _0383_ VPWR VGND sg13g2_a21o_1
X_4573_ net1155 net1068 _0320_ VPWR VGND sg13g2_nor2b_1
X_3524_ net1313 VPWR _1943_ VGND _1940_ _1942_ sg13g2_o21ai_1
X_3455_ VGND VPWR _1787_ _1876_ _1877_ net994 sg13g2_a21oi_1
X_3386_ net994 VPWR _1817_ VGND net1226 net984 sg13g2_o21ai_1
X_6174_ net98 VGND VPWR net320 s0.was_valid_out\[3\][0] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5125_ VPWR _0093_ _0819_ VGND sg13g2_inv_1
X_5056_ VGND VPWR _0761_ net1209 net299 sg13g2_or2_1
X_4007_ s0.data_out\[1\]\[4\] s0.data_out\[0\]\[4\] net948 _2380_ VPWR VGND sg13g2_mux2_1
XFILLER_25_345 VPWR VGND sg13g2_fill_1
XFILLER_13_529 VPWR VGND sg13g2_fill_2
X_5958_ net59 VGND VPWR net362 s0.data_out\[21\]\[5\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_4909_ _0571_ _0624_ net1250 _0626_ VPWR VGND sg13g2_nand3_1
X_5889_ net1016 s0.data_out\[7\]\[4\] _1507_ VPWR VGND sg13g2_and2_1
XFILLER_21_551 VPWR VGND sg13g2_fill_1
XFILLER_21_562 VPWR VGND sg13g2_decap_4
XFILLER_4_205 VPWR VGND sg13g2_fill_2
XFILLER_20_10 VPWR VGND sg13g2_decap_4
XFILLER_0_400 VPWR VGND sg13g2_decap_4
XFILLER_49_905 VPWR VGND sg13g2_decap_8
XFILLER_1_956 VPWR VGND sg13g2_decap_8
XFILLER_48_415 VPWR VGND sg13g2_decap_8
Xhold30 s0.was_valid_out\[7\][0] VPWR VGND net326 sg13g2_dlygate4sd3_1
XFILLER_0_466 VPWR VGND sg13g2_decap_8
Xhold41 s0.valid_out\[19\][0] VPWR VGND net337 sg13g2_dlygate4sd3_1
XFILLER_29_41 VPWR VGND sg13g2_fill_2
Xhold74 s0.data_out\[21\]\[1\] VPWR VGND net370 sg13g2_dlygate4sd3_1
XFILLER_21_1011 VPWR VGND sg13g2_decap_8
Xhold63 s0.data_out\[21\]\[4\] VPWR VGND net359 sg13g2_dlygate4sd3_1
Xhold52 s0.data_out\[0\]\[3\] VPWR VGND net348 sg13g2_dlygate4sd3_1
Xhold85 s0.was_valid_out\[15\][0] VPWR VGND net381 sg13g2_dlygate4sd3_1
Xhold96 s0.data_out\[0\]\[1\] VPWR VGND net392 sg13g2_dlygate4sd3_1
XFILLER_16_323 VPWR VGND sg13g2_fill_2
XFILLER_17_824 VPWR VGND sg13g2_fill_1
XFILLER_17_846 VPWR VGND sg13g2_fill_1
XFILLER_45_84 VPWR VGND sg13g2_decap_8
XFILLER_43_153 VPWR VGND sg13g2_decap_8
XFILLER_8_522 VPWR VGND sg13g2_decap_8
XFILLER_6_23 VPWR VGND sg13g2_fill_2
XFILLER_4_761 VPWR VGND sg13g2_decap_8
X_6075__204 VPWR VGND net204 sg13g2_tiehi
X_3240_ _1684_ net1006 _1645_ _1685_ VPWR VGND sg13g2_a21o_1
XFILLER_39_404 VPWR VGND sg13g2_decap_8
XFILLER_20_4 VPWR VGND sg13g2_fill_2
X_3171_ _1620_ VPWR _1621_ VGND _1616_ _1619_ sg13g2_o21ai_1
Xfanout1050 net1052 net1050 VPWR VGND sg13g2_buf_8
Xfanout1072 net605 net1072 VPWR VGND sg13g2_buf_8
Xfanout1061 net1064 net1061 VPWR VGND sg13g2_buf_8
Xfanout1083 net358 net1083 VPWR VGND sg13g2_buf_8
Xfanout1094 net1095 net1094 VPWR VGND sg13g2_buf_2
XFILLER_35_632 VPWR VGND sg13g2_fill_2
XFILLER_19_183 VPWR VGND sg13g2_fill_1
X_5812_ _1437_ net1028 _1409_ _1438_ VPWR VGND sg13g2_a21o_1
XFILLER_23_849 VPWR VGND sg13g2_decap_8
X_5743_ net1030 net1067 _1375_ VPWR VGND sg13g2_nor2b_1
X_5674_ s0.data_out\[10\]\[6\] s0.data_out\[9\]\[6\] net1043 _1319_ VPWR VGND sg13g2_mux2_1
X_4625_ _0365_ VPWR _0366_ VGND net1163 _2484_ sg13g2_o21ai_1
X_4556_ _0305_ net925 _0304_ VPWR VGND sg13g2_nand2_1
X_3507_ _1928_ _1902_ _1927_ VPWR VGND sg13g2_nand2_1
X_4487_ VPWR _0034_ net575 VGND sg13g2_inv_1
XFILLER_44_1011 VPWR VGND sg13g2_decap_8
X_3438_ s0.data_out\[4\]\[5\] s0.data_out\[5\]\[5\] net998 _1862_ VPWR VGND sg13g2_mux2_1
X_6157_ net116 VGND VPWR _0207_ s0.data_out\[5\]\[5\] clknet_leaf_13_clk sg13g2_dfrbpq_2
X_3369_ _1802_ net1250 _1801_ VPWR VGND sg13g2_nand2_1
XFILLER_46_908 VPWR VGND sg13g2_decap_8
X_5108_ _0804_ VPWR _0805_ VGND _0800_ _0803_ sg13g2_o21ai_1
X_6088_ net190 VGND VPWR _0138_ s0.data_out\[10\]\[3\] clknet_leaf_21_clk sg13g2_dfrbpq_2
XFILLER_39_993 VPWR VGND sg13g2_decap_8
X_5039_ VGND VPWR net1126 _0743_ _0744_ _0682_ sg13g2_a21oi_1
XFILLER_26_654 VPWR VGND sg13g2_fill_2
XFILLER_15_65 VPWR VGND sg13g2_fill_2
XFILLER_22_882 VPWR VGND sg13g2_fill_1
XFILLER_21_392 VPWR VGND sg13g2_fill_1
XFILLER_31_64 VPWR VGND sg13g2_decap_8
Xoutput7 net7 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_1_753 VPWR VGND sg13g2_decap_8
XFILLER_49_702 VPWR VGND sg13g2_decap_8
XFILLER_0_296 VPWR VGND sg13g2_fill_1
XFILLER_49_779 VPWR VGND sg13g2_decap_8
XFILLER_36_418 VPWR VGND sg13g2_decap_4
XFILLER_45_963 VPWR VGND sg13g2_decap_8
X_5986__29 VPWR VGND net29 sg13g2_tiehi
XFILLER_29_492 VPWR VGND sg13g2_decap_8
XFILLER_16_164 VPWR VGND sg13g2_decap_8
XFILLER_16_175 VPWR VGND sg13g2_fill_2
XFILLER_16_186 VPWR VGND sg13g2_fill_2
XFILLER_13_860 VPWR VGND sg13g2_fill_2
XFILLER_32_668 VPWR VGND sg13g2_fill_1
X_4410_ VGND VPWR _2738_ net1208 net301 sg13g2_or2_1
X_5390_ VGND VPWR _1060_ net594 net1336 sg13g2_or2_1
X_4341_ net1196 VPWR _2672_ VGND _2670_ _2671_ sg13g2_o21ai_1
X_4272_ net1260 _2587_ _2612_ VPWR VGND sg13g2_nor2_1
XFILLER_28_1028 VPWR VGND sg13g2_fill_1
X_6011_ net274 VGND VPWR net322 s0.was_valid_out\[16\][0] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_3223_ _1668_ net1264 _1667_ VPWR VGND sg13g2_nand2_1
X_3154_ _1602_ _1605_ net1327 _1606_ VPWR VGND sg13g2_nand3_1
XFILLER_36_952 VPWR VGND sg13g2_decap_8
XFILLER_22_167 VPWR VGND sg13g2_fill_1
X_3987_ VPWR VGND _2358_ _2359_ _2354_ net1211 _2360_ _2350_ sg13g2_a221oi_1
X_5726_ net1023 s0.data_out\[8\]\[0\] _1360_ VPWR VGND sg13g2_and2_1
X_5657_ _1247_ _1301_ _1302_ VPWR VGND sg13g2_and2_1
XFILLER_2_506 VPWR VGND sg13g2_decap_4
X_4608_ VGND VPWR _0351_ net558 net1302 sg13g2_or2_1
X_5588_ net1035 s0.data_out\[9\]\[0\] _1241_ VPWR VGND sg13g2_and2_1
X_4539_ _0292_ _2742_ _0290_ _0291_ VPWR VGND sg13g2_and3_1
X_6209_ net247 VGND VPWR _0259_ s0.genblk1\[19\].modules.bubble clknet_leaf_3_clk
+ sg13g2_dfrbpq_1
XFILLER_46_705 VPWR VGND sg13g2_decap_8
XFILLER_26_42 VPWR VGND sg13g2_decap_8
XFILLER_42_922 VPWR VGND sg13g2_decap_8
Xclkbuf_3_6__f_clk clknet_0_clk clknet_3_6__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_41_410 VPWR VGND sg13g2_fill_1
XFILLER_26_86 VPWR VGND sg13g2_decap_8
XFILLER_26_495 VPWR VGND sg13g2_decap_8
XFILLER_42_999 VPWR VGND sg13g2_decap_8
XFILLER_42_85 VPWR VGND sg13g2_fill_1
XFILLER_6_845 VPWR VGND sg13g2_fill_2
XFILLER_6_834 VPWR VGND sg13g2_decap_8
X_6072__207 VPWR VGND net207 sg13g2_tiehi
XFILLER_1_550 VPWR VGND sg13g2_decap_8
XFILLER_3_79 VPWR VGND sg13g2_fill_2
XFILLER_49_576 VPWR VGND sg13g2_decap_8
XFILLER_45_760 VPWR VGND sg13g2_decap_8
XFILLER_17_451 VPWR VGND sg13g2_decap_8
XFILLER_33_900 VPWR VGND sg13g2_decap_4
XFILLER_44_270 VPWR VGND sg13g2_decap_8
X_4890_ VGND VPWR net1149 _0606_ _0607_ _0557_ sg13g2_a21oi_1
X_3910_ s0.data_out\[0\]\[0\] s0.data_out\[1\]\[0\] net955 _2291_ VPWR VGND sg13g2_mux2_1
X_3841_ net953 net1045 _2227_ VPWR VGND sg13g2_nor2b_1
X_3772_ _2167_ net1222 net956 VPWR VGND sg13g2_nand2_1
XFILLER_32_476 VPWR VGND sg13g2_decap_8
X_5511_ VGND VPWR net1081 net521 _1170_ _1169_ sg13g2_a21oi_1
X_5442_ VGND VPWR _1104_ _1110_ _1111_ _1094_ sg13g2_a21oi_1
X_5373_ net1339 VPWR _1045_ VGND net938 _1044_ sg13g2_o21ai_1
X_4324_ VGND VPWR net1179 s0.data_out\[19\]\[3\] _2657_ _2656_ sg13g2_a21oi_1
XFILLER_41_1003 VPWR VGND sg13g2_decap_8
X_4255_ _2595_ net1200 net592 VPWR VGND sg13g2_nand2_1
X_4186_ _2531_ VPWR _2532_ VGND net1206 s0.data_out\[20\]\[2\] sg13g2_o21ai_1
X_3206_ _1650_ VPWR _1651_ VGND net1008 _2491_ sg13g2_o21ai_1
XFILLER_28_705 VPWR VGND sg13g2_decap_8
X_3137_ _1586_ _1591_ _1592_ VPWR VGND sg13g2_nor2_1
XFILLER_27_237 VPWR VGND sg13g2_fill_2
X_5973__43 VPWR VGND net43 sg13g2_tiehi
XFILLER_23_487 VPWR VGND sg13g2_decap_8
X_5709_ net1223 net1049 _1347_ VPWR VGND sg13g2_nor2_1
XFILLER_12_88 VPWR VGND sg13g2_fill_2
XFILLER_3_859 VPWR VGND sg13g2_decap_8
Xhold160 s0.data_out\[16\]\[5\] VPWR VGND net456 sg13g2_dlygate4sd3_1
Xhold171 s0.data_out\[7\]\[2\] VPWR VGND net467 sg13g2_dlygate4sd3_1
Xhold182 s0.data_out\[18\]\[3\] VPWR VGND net478 sg13g2_dlygate4sd3_1
Xhold193 _2196_ VPWR VGND net489 sg13g2_dlygate4sd3_1
XFILLER_19_727 VPWR VGND sg13g2_fill_1
XFILLER_46_557 VPWR VGND sg13g2_fill_1
XFILLER_46_546 VPWR VGND sg13g2_decap_8
XFILLER_27_760 VPWR VGND sg13g2_fill_2
XFILLER_26_270 VPWR VGND sg13g2_decap_8
XFILLER_41_240 VPWR VGND sg13g2_fill_1
XFILLER_30_947 VPWR VGND sg13g2_fill_1
XFILLER_10_693 VPWR VGND sg13g2_fill_2
X_4040_ _2407_ net940 net1065 VPWR VGND sg13g2_nand2_1
XFILLER_49_373 VPWR VGND sg13g2_decap_8
X_5991_ net23 VGND VPWR _0041_ s0.data_out\[18\]\[2\] clknet_leaf_35_clk sg13g2_dfrbpq_2
X_4942_ net1138 VPWR _0655_ VGND _0653_ _0654_ sg13g2_o21ai_1
X_4873_ VPWR _0070_ _0590_ VGND sg13g2_inv_1
X_3824_ _2212_ net930 _2211_ VPWR VGND sg13g2_nand2_1
X_6124__152 VPWR VGND net152 sg13g2_tiehi
X_3755_ s0.data_out\[3\]\[5\] s0.data_out\[2\]\[5\] net966 _2152_ VPWR VGND sg13g2_mux2_1
X_5970__46 VPWR VGND net46 sg13g2_tiehi
X_3686_ _2087_ VPWR _2088_ VGND _2083_ _2086_ sg13g2_o21ai_1
X_5425_ _1091_ _1092_ _1094_ VPWR VGND _1093_ sg13g2_nand3b_1
X_5356_ net1089 net1062 _1030_ VPWR VGND sg13g2_nor2b_1
X_4307_ net1178 s0.data_out\[19\]\[1\] _2642_ VPWR VGND sg13g2_and2_1
X_5287_ VGND VPWR net1117 _0967_ _0968_ _0938_ sg13g2_a21oi_1
X_4238_ s0.data_out\[21\]\[0\] s0.data_out\[20\]\[0\] net1198 _2578_ VPWR VGND sg13g2_mux2_1
X_4169_ net368 net1206 _2517_ VPWR VGND sg13g2_nor2b_1
XFILLER_16_708 VPWR VGND sg13g2_decap_8
XFILLER_24_752 VPWR VGND sg13g2_fill_2
XFILLER_12_936 VPWR VGND sg13g2_decap_8
XFILLER_23_262 VPWR VGND sg13g2_decap_4
XFILLER_8_929 VPWR VGND sg13g2_decap_8
XFILLER_47_822 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_19_546 VPWR VGND sg13g2_fill_2
XFILLER_47_899 VPWR VGND sg13g2_decap_8
XFILLER_0_69 VPWR VGND sg13g2_decap_4
XFILLER_0_47 VPWR VGND sg13g2_decap_4
XFILLER_46_398 VPWR VGND sg13g2_decap_8
XFILLER_15_752 VPWR VGND sg13g2_decap_4
XFILLER_15_774 VPWR VGND sg13g2_fill_1
XFILLER_15_785 VPWR VGND sg13g2_decap_4
X_6108__169 VPWR VGND net169 sg13g2_tiehi
XFILLER_14_284 VPWR VGND sg13g2_fill_2
XFILLER_30_744 VPWR VGND sg13g2_decap_4
XFILLER_31_1013 VPWR VGND sg13g2_decap_8
X_3540_ _1952_ _1955_ net1312 _1956_ VPWR VGND sg13g2_nand3_1
X_5210_ net1100 net1070 _0898_ VPWR VGND sg13g2_nor2b_1
XFILLER_6_494 VPWR VGND sg13g2_fill_2
X_3471_ s0.data_out\[5\]\[0\] s0.data_out\[4\]\[0\] net989 _1892_ VPWR VGND sg13g2_mux2_1
X_6190_ net80 VGND VPWR _0240_ s0.data_out\[2\]\[2\] clknet_leaf_6_clk sg13g2_dfrbpq_2
X_5141_ s0.data_out\[14\]\[0\] s0.data_out\[13\]\[0\] net1119 _0834_ VPWR VGND sg13g2_mux2_1
X_5072_ net1113 s0.data_out\[13\]\[0\] _0773_ VPWR VGND sg13g2_and2_1
X_4023_ VPWR VGND _2379_ _2395_ _2394_ _2368_ _2396_ _2393_ sg13g2_a221oi_1
XFILLER_38_899 VPWR VGND sg13g2_fill_1
XFILLER_37_343 VPWR VGND sg13g2_decap_8
XFILLER_25_538 VPWR VGND sg13g2_decap_4
X_5974_ net42 VGND VPWR _0024_ s0.genblk1\[1\].modules.bubble clknet_leaf_10_clk sg13g2_dfrbpq_1
X_4925_ net1319 net299 _0072_ VPWR VGND sg13g2_and2_1
XFILLER_20_221 VPWR VGND sg13g2_decap_8
X_4856_ _0575_ VPWR _0576_ VGND net1323 net456 sg13g2_o21ai_1
XFILLER_21_777 VPWR VGND sg13g2_decap_8
XFILLER_21_788 VPWR VGND sg13g2_fill_1
XFILLER_21_799 VPWR VGND sg13g2_fill_1
X_3807_ s0.data_out\[1\]\[3\] s0.data_out\[2\]\[3\] net965 _2197_ VPWR VGND sg13g2_mux2_1
X_4787_ net1248 _0514_ _0516_ VPWR VGND sg13g2_nor2_1
X_3738_ _2134_ VPWR _2135_ VGND net1211 _2120_ sg13g2_o21ai_1
X_3669_ _2069_ _2072_ net1307 _2073_ VPWR VGND sg13g2_nand3_1
X_5408_ _1077_ net1096 net486 VPWR VGND sg13g2_nand2_1
X_5339_ net1088 net1070 _1015_ VPWR VGND sg13g2_nor2b_1
XFILLER_48_619 VPWR VGND sg13g2_decap_8
XFILLER_28_321 VPWR VGND sg13g2_fill_2
XFILLER_29_855 VPWR VGND sg13g2_decap_8
XFILLER_29_888 VPWR VGND sg13g2_fill_1
XFILLER_44_836 VPWR VGND sg13g2_decap_8
XFILLER_43_357 VPWR VGND sg13g2_decap_4
XFILLER_15_1008 VPWR VGND sg13g2_decap_8
XFILLER_11_265 VPWR VGND sg13g2_decap_8
XFILLER_7_258 VPWR VGND sg13g2_decap_8
XFILLER_4_921 VPWR VGND sg13g2_decap_8
XFILLER_4_998 VPWR VGND sg13g2_decap_8
Xfanout1232 net1234 net1232 VPWR VGND sg13g2_buf_2
Xfanout1221 _2450_ net1221 VPWR VGND sg13g2_buf_8
Xfanout1210 _2621_ net1210 VPWR VGND sg13g2_buf_8
Xfanout1243 net1245 net1243 VPWR VGND sg13g2_buf_8
Xfanout1254 net1259 net1254 VPWR VGND sg13g2_buf_8
Xfanout1265 net1267 net1265 VPWR VGND sg13g2_buf_8
Xfanout1298 net1299 net1298 VPWR VGND sg13g2_buf_8
Xfanout1287 net1288 net1287 VPWR VGND sg13g2_buf_8
Xfanout1276 ui_in[1] net1276 VPWR VGND sg13g2_buf_8
XFILLER_47_696 VPWR VGND sg13g2_decap_8
XFILLER_15_571 VPWR VGND sg13g2_decap_8
XFILLER_43_891 VPWR VGND sg13g2_decap_8
X_4710_ net922 _2485_ _0444_ VPWR VGND sg13g2_nor2_1
X_5690_ _1275_ _1334_ net1252 _1335_ VPWR VGND sg13g2_nand3_1
X_4641_ s0.data_out\[18\]\[7\] s0.data_out\[17\]\[7\] net1163 _0382_ VPWR VGND sg13g2_mux2_1
X_6121__155 VPWR VGND net155 sg13g2_tiehi
X_4572_ VGND VPWR _2804_ _0318_ _0319_ net1169 sg13g2_a21oi_1
X_3523_ _1941_ VPWR _1942_ VGND _1936_ _1939_ sg13g2_o21ai_1
X_3454_ _1876_ net535 net998 VPWR VGND sg13g2_nand2b_1
XFILLER_6_291 VPWR VGND sg13g2_decap_8
XFILLER_41_0 VPWR VGND sg13g2_fill_2
X_3385_ net1313 net318 _0199_ VPWR VGND sg13g2_and2_1
X_6173_ net99 VGND VPWR _0223_ s0.genblk1\[3\].modules.bubble clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5124_ _0818_ VPWR _0819_ VGND _0814_ _0817_ sg13g2_o21ai_1
X_5055_ _0645_ _0758_ _0759_ _0760_ VPWR VGND sg13g2_nor3_1
X_4006_ _2379_ _2375_ _2376_ _2377_ VPWR VGND sg13g2_and3_1
XFILLER_37_184 VPWR VGND sg13g2_decap_8
XFILLER_13_508 VPWR VGND sg13g2_decap_8
X_5957_ net60 VGND VPWR net360 s0.data_out\[21\]\[4\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_4908_ VGND VPWR _0571_ _0624_ _0625_ net1250 sg13g2_a21oi_1
X_5888_ _1506_ _2467_ _1505_ VPWR VGND sg13g2_nand2_1
X_4839_ _0561_ net1220 _2485_ VPWR VGND sg13g2_nand2_1
X_6509_ s0.was_valid_out\[21\][0] net1 VPWR VGND sg13g2_buf_1
XFILLER_1_935 VPWR VGND sg13g2_decap_8
XFILLER_0_445 VPWR VGND sg13g2_decap_8
Xhold31 _0176_ VPWR VGND net327 sg13g2_dlygate4sd3_1
Xhold20 s0.genblk1\[11\].modules.bubble VPWR VGND net316 sg13g2_dlygate4sd3_1
XFILLER_29_31 VPWR VGND sg13g2_fill_1
Xhold53 s0.data_out\[2\]\[5\] VPWR VGND net349 sg13g2_dlygate4sd3_1
Xhold42 s0.shift_out\[16\][0] VPWR VGND net338 sg13g2_dlygate4sd3_1
Xhold64 _0007_ VPWR VGND net360 sg13g2_dlygate4sd3_1
Xhold97 s0.was_valid_out\[2\][0] VPWR VGND net393 sg13g2_dlygate4sd3_1
Xhold75 _2527_ VPWR VGND net371 sg13g2_dlygate4sd3_1
Xhold86 _0073_ VPWR VGND net382 sg13g2_dlygate4sd3_1
XFILLER_45_30 VPWR VGND sg13g2_fill_2
X_6068__212 VPWR VGND net212 sg13g2_tiehi
XFILLER_44_655 VPWR VGND sg13g2_decap_8
XFILLER_43_143 VPWR VGND sg13g2_decap_4
XFILLER_16_346 VPWR VGND sg13g2_fill_2
XFILLER_17_869 VPWR VGND sg13g2_decap_8
XFILLER_8_589 VPWR VGND sg13g2_fill_1
XFILLER_8_567 VPWR VGND sg13g2_fill_1
XFILLER_39_416 VPWR VGND sg13g2_decap_8
XFILLER_6_1028 VPWR VGND sg13g2_fill_1
XFILLER_6_1017 VPWR VGND sg13g2_decap_8
X_3170_ VGND VPWR _1620_ net503 net1327 sg13g2_or2_1
Xfanout1040 s0.shift_out\[9\][0] net1040 VPWR VGND sg13g2_buf_8
Xfanout1051 net1052 net1051 VPWR VGND sg13g2_buf_8
Xfanout1062 net1064 net1062 VPWR VGND sg13g2_buf_8
Xfanout1073 net1076 net1073 VPWR VGND sg13g2_buf_8
Xfanout1095 s0.shift_out\[11\][0] net1095 VPWR VGND sg13g2_buf_1
Xfanout1084 net1087 net1084 VPWR VGND sg13g2_buf_8
XFILLER_48_983 VPWR VGND sg13g2_decap_8
XFILLER_47_460 VPWR VGND sg13g2_fill_1
XFILLER_35_644 VPWR VGND sg13g2_fill_2
XFILLER_34_121 VPWR VGND sg13g2_decap_4
X_5811_ s0.data_out\[9\]\[7\] s0.data_out\[8\]\[7\] net1032 _1437_ VPWR VGND sg13g2_mux2_1
X_5742_ net1024 net608 _1374_ VPWR VGND sg13g2_and2_1
XFILLER_34_198 VPWR VGND sg13g2_fill_1
X_5673_ _1318_ net1041 net542 VPWR VGND sg13g2_nand2_1
X_4624_ _0365_ net1163 net496 VPWR VGND sg13g2_nand2_1
X_4555_ s0.data_out\[17\]\[0\] s0.data_out\[18\]\[0\] net1175 _0304_ VPWR VGND sg13g2_mux2_1
X_3506_ _1914_ _1923_ _1924_ _1926_ _1927_ VPWR VGND sg13g2_nor4_1
X_4486_ _2802_ VPWR _2803_ VGND _2798_ _2801_ sg13g2_o21ai_1
X_3437_ VPWR _0206_ _1861_ VGND sg13g2_inv_1
X_3368_ VGND VPWR net1004 _1800_ _1801_ _1748_ sg13g2_a21oi_1
X_6156_ net117 VGND VPWR _0206_ s0.data_out\[5\]\[4\] clknet_leaf_14_clk sg13g2_dfrbpq_2
X_5107_ VGND VPWR _0804_ net525 net1322 sg13g2_or2_1
X_6210__234 VPWR VGND net234 sg13g2_tiehi
XFILLER_39_972 VPWR VGND sg13g2_decap_8
X_6087_ net191 VGND VPWR _0137_ s0.data_out\[10\]\[2\] clknet_leaf_21_clk sg13g2_dfrbpq_2
X_3299_ net1000 VPWR _1737_ VGND _1735_ _1736_ sg13g2_o21ai_1
XFILLER_38_482 VPWR VGND sg13g2_fill_2
X_5038_ s0.data_out\[15\]\[4\] s0.data_out\[14\]\[4\] net1133 _0743_ VPWR VGND sg13g2_mux2_1
XFILLER_38_493 VPWR VGND sg13g2_fill_1
XFILLER_25_132 VPWR VGND sg13g2_decap_8
XFILLER_26_688 VPWR VGND sg13g2_fill_2
XFILLER_40_135 VPWR VGND sg13g2_fill_2
XFILLER_40_102 VPWR VGND sg13g2_fill_2
XFILLER_31_32 VPWR VGND sg13g2_fill_1
Xoutput8 net8 uo_out[6] VPWR VGND sg13g2_buf_1
XFILLER_1_732 VPWR VGND sg13g2_decap_8
XFILLER_0_253 VPWR VGND sg13g2_decap_8
XFILLER_49_758 VPWR VGND sg13g2_decap_8
XFILLER_45_942 VPWR VGND sg13g2_decap_8
XFILLER_17_633 VPWR VGND sg13g2_decap_4
XFILLER_16_143 VPWR VGND sg13g2_decap_8
XFILLER_44_485 VPWR VGND sg13g2_fill_2
XFILLER_16_198 VPWR VGND sg13g2_decap_4
XFILLER_32_647 VPWR VGND sg13g2_decap_8
XFILLER_12_393 VPWR VGND sg13g2_fill_2
X_4340_ net1182 net1053 _2671_ VPWR VGND sg13g2_nor2b_1
XFILLER_28_1007 VPWR VGND sg13g2_decap_8
XFILLER_4_592 VPWR VGND sg13g2_decap_4
X_4271_ _2611_ _2606_ _2610_ VPWR VGND sg13g2_nand2_1
X_6010_ net275 VGND VPWR _0060_ s0.genblk1\[16\].modules.bubble clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
X_3222_ VGND VPWR net1014 _1666_ _1667_ _1616_ sg13g2_a21oi_1
X_3153_ net1012 VPWR _1605_ VGND _1603_ _1604_ sg13g2_o21ai_1
XFILLER_28_909 VPWR VGND sg13g2_decap_8
XFILLER_48_780 VPWR VGND sg13g2_decap_8
XFILLER_35_463 VPWR VGND sg13g2_decap_8
X_5985__30 VPWR VGND net30 sg13g2_tiehi
XFILLER_23_669 VPWR VGND sg13g2_decap_4
X_3986_ VGND VPWR _2299_ _2353_ _2359_ net1274 sg13g2_a21oi_1
X_5725_ _1359_ net919 _1358_ VPWR VGND sg13g2_nand2_1
X_5656_ _1301_ net1078 _1300_ VPWR VGND sg13g2_nand2b_1
X_4607_ net1301 VPWR _0350_ VGND _2461_ _0349_ sg13g2_o21ai_1
X_5587_ _1240_ net934 _1239_ VPWR VGND sg13g2_nand2_1
X_4538_ _0291_ _0272_ _2833_ VPWR VGND sg13g2_nand2b_1
X_4469_ VGND VPWR _2788_ net586 net1290 sg13g2_or2_1
X_6208_ net260 VGND VPWR _0258_ s0.shift_out\[1\][0] clknet_leaf_10_clk sg13g2_dfrbpq_2
X_6139_ net135 VGND VPWR _0189_ s0.valid_out\[6\][0] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_42_901 VPWR VGND sg13g2_decap_8
XFILLER_26_441 VPWR VGND sg13g2_decap_8
X_6065__215 VPWR VGND net215 sg13g2_tiehi
XFILLER_42_978 VPWR VGND sg13g2_decap_8
XFILLER_42_20 VPWR VGND sg13g2_decap_4
XFILLER_41_455 VPWR VGND sg13g2_fill_1
XFILLER_41_477 VPWR VGND sg13g2_decap_4
XFILLER_10_831 VPWR VGND sg13g2_decap_8
XFILLER_5_378 VPWR VGND sg13g2_fill_2
XFILLER_3_25 VPWR VGND sg13g2_fill_2
XFILLER_3_14 VPWR VGND sg13g2_fill_2
XFILLER_49_555 VPWR VGND sg13g2_decap_8
XFILLER_17_496 VPWR VGND sg13g2_decap_4
X_3840_ VGND VPWR _2136_ _2225_ _2226_ net962 sg13g2_a21oi_1
XFILLER_32_455 VPWR VGND sg13g2_fill_2
X_3771_ net962 VPWR _2166_ VGND net1225 net953 sg13g2_o21ai_1
X_5982__33 VPWR VGND net33 sg13g2_tiehi
X_5510_ net1081 net1051 _1169_ VPWR VGND sg13g2_nor2b_1
X_5441_ _1110_ _1105_ _1099_ VPWR VGND sg13g2_nand2b_1
X_5372_ VGND VPWR net1091 s0.data_out\[11\]\[5\] _1044_ _1043_ sg13g2_a21oi_1
X_4323_ net1179 net1061 _2656_ VPWR VGND sg13g2_nor2b_1
X_4254_ VGND VPWR net1203 _2593_ _2594_ _2568_ sg13g2_a21oi_1
X_4185_ VGND VPWR net1206 _2479_ _2531_ net1203 sg13g2_a21oi_1
X_3205_ _1650_ net1011 net484 VPWR VGND sg13g2_nand2_1
X_3136_ VGND VPWR net1222 net1020 _1591_ net1015 sg13g2_a21oi_1
XFILLER_24_923 VPWR VGND sg13g2_fill_2
XFILLER_11_606 VPWR VGND sg13g2_decap_4
XFILLER_23_466 VPWR VGND sg13g2_fill_1
X_3969_ VGND VPWR net945 net334 _2343_ _2342_ sg13g2_a21oi_1
X_5708_ net1053 net1246 net1223 _0149_ VPWR VGND sg13g2_mux2_1
X_5639_ VGND VPWR _1286_ net521 net1346 sg13g2_or2_1
XFILLER_12_56 VPWR VGND sg13g2_fill_2
XFILLER_3_838 VPWR VGND sg13g2_decap_8
Xhold161 s0.data_out\[14\]\[0\] VPWR VGND net457 sg13g2_dlygate4sd3_1
Xhold150 s0.data_out\[2\]\[3\] VPWR VGND net446 sg13g2_dlygate4sd3_1
Xhold183 s0.data_out\[1\]\[5\] VPWR VGND net479 sg13g2_dlygate4sd3_1
Xhold194 s0.data_out\[20\]\[2\] VPWR VGND net490 sg13g2_dlygate4sd3_1
Xhold172 s0.data_out\[17\]\[0\] VPWR VGND net468 sg13g2_dlygate4sd3_1
XFILLER_18_249 VPWR VGND sg13g2_fill_1
XFILLER_14_433 VPWR VGND sg13g2_fill_2
XFILLER_6_632 VPWR VGND sg13g2_decap_4
XFILLER_45_7 VPWR VGND sg13g2_fill_1
XFILLER_2_882 VPWR VGND sg13g2_decap_8
XFILLER_37_514 VPWR VGND sg13g2_decap_4
XFILLER_37_558 VPWR VGND sg13g2_decap_8
X_5990_ net24 VGND VPWR _0040_ s0.data_out\[18\]\[1\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_4941_ net1122 net1074 _0654_ VPWR VGND sg13g2_nor2b_1
XFILLER_17_260 VPWR VGND sg13g2_fill_2
X_4872_ _0589_ VPWR _0590_ VGND _0585_ _0588_ sg13g2_o21ai_1
X_3823_ s0.data_out\[1\]\[5\] s0.data_out\[2\]\[5\] net966 _2211_ VPWR VGND sg13g2_mux2_1
X_3754_ _2090_ _2150_ _2151_ VPWR VGND sg13g2_and2_1
X_3685_ VGND VPWR _2087_ net509 net1308 sg13g2_or2_1
X_5424_ net1242 _1090_ _1093_ VPWR VGND sg13g2_nor2_1
X_5355_ net1088 net613 _1029_ VPWR VGND sg13g2_and2_1
X_4306_ _2641_ net931 _2640_ VPWR VGND sg13g2_nand2_1
X_5286_ _0966_ net1107 _0939_ _0967_ VPWR VGND sg13g2_a21o_1
X_4237_ _2525_ _2576_ net1273 _2577_ VPWR VGND sg13g2_nand3_1
X_4168_ net1202 VPWR _2516_ VGND _2514_ _2515_ sg13g2_o21ai_1
XFILLER_28_558 VPWR VGND sg13g2_decap_8
X_4099_ _2458_ net962 VPWR VGND sg13g2_inv_2
X_3119_ _1573_ VPWR _1576_ VGND net1266 _1549_ sg13g2_o21ai_1
XFILLER_24_742 VPWR VGND sg13g2_fill_2
X_6062__218 VPWR VGND net218 sg13g2_tiehi
XFILLER_3_613 VPWR VGND sg13g2_decap_4
XFILLER_3_679 VPWR VGND sg13g2_fill_2
XFILLER_24_1021 VPWR VGND sg13g2_decap_8
XFILLER_47_801 VPWR VGND sg13g2_decap_8
XFILLER_47_878 VPWR VGND sg13g2_decap_8
XFILLER_11_981 VPWR VGND sg13g2_decap_8
XFILLER_7_985 VPWR VGND sg13g2_decap_8
X_3470_ _1835_ _1890_ _1891_ VPWR VGND sg13g2_and2_1
X_5140_ VGND VPWR net1127 _0832_ _0833_ _0779_ sg13g2_a21oi_1
X_5071_ _0772_ net937 _0771_ VPWR VGND sg13g2_nand2_1
XFILLER_29_2 VPWR VGND sg13g2_fill_1
X_4022_ _2285_ VPWR _2395_ VGND _2375_ _2378_ sg13g2_o21ai_1
XFILLER_49_182 VPWR VGND sg13g2_decap_8
XFILLER_49_160 VPWR VGND sg13g2_decap_8
XFILLER_37_311 VPWR VGND sg13g2_fill_1
X_5973_ net43 VGND VPWR _0023_ s0.shift_out\[20\][0] clknet_leaf_1_clk sg13g2_dfrbpq_2
X_4924_ VGND VPWR _0635_ _0639_ _0071_ _0640_ sg13g2_a21oi_1
X_4855_ _0571_ _0574_ net1323 _0575_ VPWR VGND sg13g2_nand3_1
X_4786_ _0515_ net1248 _0514_ VPWR VGND sg13g2_nand2_1
XFILLER_20_266 VPWR VGND sg13g2_fill_2
X_3806_ VPWR _0240_ net489 VGND sg13g2_inv_1
X_3737_ _2134_ net1262 _2133_ VPWR VGND sg13g2_nand2_1
X_3668_ net971 VPWR _2072_ VGND _2070_ _2071_ sg13g2_o21ai_1
X_5407_ _1066_ _1074_ _1075_ _1076_ VPWR VGND sg13g2_nor3_1
X_3599_ s0.data_out\[4\]\[0\] s0.data_out\[3\]\[0\] net976 _2008_ VPWR VGND sg13g2_mux2_1
X_5338_ VGND VPWR _0948_ _1013_ _1014_ net1102 sg13g2_a21oi_1
XFILLER_0_649 VPWR VGND sg13g2_decap_8
X_5269_ VGND VPWR net1100 _0949_ _0950_ _0898_ sg13g2_a21oi_1
XFILLER_18_33 VPWR VGND sg13g2_fill_1
XFILLER_44_815 VPWR VGND sg13g2_decap_8
XFILLER_16_506 VPWR VGND sg13g2_fill_2
XFILLER_43_314 VPWR VGND sg13g2_decap_8
XFILLER_16_517 VPWR VGND sg13g2_decap_8
XFILLER_34_65 VPWR VGND sg13g2_decap_8
X_6107__170 VPWR VGND net170 sg13g2_tiehi
XFILLER_7_215 VPWR VGND sg13g2_decap_4
XFILLER_4_900 VPWR VGND sg13g2_decap_8
XFILLER_3_421 VPWR VGND sg13g2_fill_1
XFILLER_3_410 VPWR VGND sg13g2_decap_8
X_6218__110 VPWR VGND net110 sg13g2_tiehi
XFILLER_4_977 VPWR VGND sg13g2_decap_8
Xfanout1222 _2449_ net1222 VPWR VGND sg13g2_buf_8
Xfanout1211 net1212 net1211 VPWR VGND sg13g2_buf_8
Xfanout1200 net1201 net1200 VPWR VGND sg13g2_buf_8
Xfanout1233 net1234 net1233 VPWR VGND sg13g2_buf_8
Xfanout1244 net1245 net1244 VPWR VGND sg13g2_buf_8
Xfanout1255 net1259 net1255 VPWR VGND sg13g2_buf_1
Xfanout1299 net1300 net1299 VPWR VGND sg13g2_buf_8
X_6114__163 VPWR VGND net163 sg13g2_tiehi
Xfanout1288 net1290 net1288 VPWR VGND sg13g2_buf_8
Xfanout1277 net1280 net1277 VPWR VGND sg13g2_buf_8
Xfanout1266 net1267 net1266 VPWR VGND sg13g2_buf_8
XFILLER_47_675 VPWR VGND sg13g2_decap_8
XFILLER_35_859 VPWR VGND sg13g2_decap_8
XFILLER_43_870 VPWR VGND sg13g2_decap_8
XFILLER_15_594 VPWR VGND sg13g2_fill_2
X_4640_ _0381_ net1164 net341 VPWR VGND sg13g2_nand2_1
X_4571_ _0318_ s0.data_out\[17\]\[2\] net1175 VPWR VGND sg13g2_nand2b_1
X_3522_ _2471_ VPWR _1941_ VGND net319 net988 sg13g2_o21ai_1
XFILLER_7_782 VPWR VGND sg13g2_fill_2
X_3453_ VPWR _0208_ _1875_ VGND sg13g2_inv_1
X_6172_ net100 VGND VPWR _0222_ s0.shift_out\[4\][0] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_3384_ VGND VPWR _1811_ _1815_ _0198_ _1816_ sg13g2_a21oi_1
X_5123_ VGND VPWR _0818_ net598 net1321 sg13g2_or2_1
XFILLER_34_0 VPWR VGND sg13g2_decap_8
X_5054_ _0737_ _0738_ _0759_ VPWR VGND sg13g2_nor2b_1
XFILLER_29_119 VPWR VGND sg13g2_decap_8
X_4005_ VPWR _2378_ _2377_ VGND sg13g2_inv_1
XFILLER_26_804 VPWR VGND sg13g2_decap_4
XFILLER_26_859 VPWR VGND sg13g2_decap_4
XFILLER_41_829 VPWR VGND sg13g2_decap_8
XFILLER_40_306 VPWR VGND sg13g2_fill_2
X_5956_ net61 VGND VPWR net367 s0.data_out\[21\]\[3\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_5887_ s0.data_out\[7\]\[4\] s0.data_out\[8\]\[4\] net1032 _1505_ VPWR VGND sg13g2_mux2_1
X_4907_ _0624_ net1148 _0623_ VPWR VGND sg13g2_nand2b_1
X_4838_ net1317 VPWR _0560_ VGND net922 _0559_ sg13g2_o21ai_1
XFILLER_21_575 VPWR VGND sg13g2_decap_8
X_4769_ _0497_ net1146 _0465_ _0498_ VPWR VGND sg13g2_a21o_1
XFILLER_1_914 VPWR VGND sg13g2_decap_8
XFILLER_0_424 VPWR VGND sg13g2_decap_8
Xhold21 s0.genblk1\[4\].modules.bubble VPWR VGND net317 sg13g2_dlygate4sd3_1
Xhold32 s0.was_valid_out\[1\][0] VPWR VGND net328 sg13g2_dlygate4sd3_1
Xhold10 s0.genblk1\[21\].modules.bubble VPWR VGND net306 sg13g2_dlygate4sd3_1
Xhold43 s0.shift_out\[7\][0] VPWR VGND net339 sg13g2_dlygate4sd3_1
Xhold54 s0.data_out\[8\]\[4\] VPWR VGND net350 sg13g2_dlygate4sd3_1
Xhold65 s0.data_out\[21\]\[5\] VPWR VGND net361 sg13g2_dlygate4sd3_1
Xhold87 s0.was_valid_out\[5\][0] VPWR VGND net383 sg13g2_dlygate4sd3_1
Xhold98 s0.data_out\[1\]\[4\] VPWR VGND net394 sg13g2_dlygate4sd3_1
Xhold76 s0.was_valid_out\[21\][0] VPWR VGND net372 sg13g2_dlygate4sd3_1
XFILLER_17_815 VPWR VGND sg13g2_decap_8
XFILLER_16_325 VPWR VGND sg13g2_fill_1
XFILLER_16_336 VPWR VGND sg13g2_fill_1
XFILLER_16_358 VPWR VGND sg13g2_fill_1
XFILLER_8_502 VPWR VGND sg13g2_fill_2
XFILLER_8_557 VPWR VGND sg13g2_fill_2
XFILLER_3_262 VPWR VGND sg13g2_fill_1
Xfanout1030 s0.shift_out\[8\][0] net1030 VPWR VGND sg13g2_buf_8
Xfanout1041 net1044 net1041 VPWR VGND sg13g2_buf_8
Xfanout1063 net1064 net1063 VPWR VGND sg13g2_buf_8
Xfanout1074 net1076 net1074 VPWR VGND sg13g2_buf_8
Xfanout1052 net603 net1052 VPWR VGND sg13g2_buf_8
XFILLER_48_962 VPWR VGND sg13g2_decap_8
Xfanout1096 net1099 net1096 VPWR VGND sg13g2_buf_8
Xfanout1085 net1087 net1085 VPWR VGND sg13g2_buf_8
XFILLER_19_174 VPWR VGND sg13g2_decap_8
XFILLER_35_634 VPWR VGND sg13g2_fill_1
X_5810_ _1436_ net1032 net595 VPWR VGND sg13g2_nand2_1
XFILLER_35_689 VPWR VGND sg13g2_decap_8
XFILLER_34_144 VPWR VGND sg13g2_decap_8
XFILLER_34_166 VPWR VGND sg13g2_fill_2
XFILLER_37_1020 VPWR VGND sg13g2_decap_8
X_5741_ _1373_ net919 _1372_ VPWR VGND sg13g2_nand2_1
X_5672_ VGND VPWR net1083 _1316_ _1317_ _1289_ sg13g2_a21oi_1
X_4623_ VGND VPWR _0364_ _0363_ net1269 sg13g2_or2_1
X_4554_ net1219 _0298_ _0038_ VPWR VGND sg13g2_nor2_1
X_3505_ _1925_ VPWR _1926_ VGND net1267 _1900_ sg13g2_o21ai_1
X_4485_ VGND VPWR _2802_ net574 net1288 sg13g2_or2_1
X_3436_ _1860_ VPWR _1861_ VGND net1315 net402 sg13g2_o21ai_1
X_3367_ _1799_ net995 _1749_ _1800_ VPWR VGND sg13g2_a21o_1
X_6155_ net118 VGND VPWR _0205_ s0.data_out\[5\]\[3\] clknet_leaf_15_clk sg13g2_dfrbpq_2
X_5106_ net1322 VPWR _0803_ VGND _2452_ _0802_ sg13g2_o21ai_1
X_6086_ net192 VGND VPWR _0136_ s0.data_out\[10\]\[1\] clknet_leaf_21_clk sg13g2_dfrbpq_2
XFILLER_39_951 VPWR VGND sg13g2_decap_8
X_5037_ _0742_ net1132 net525 VPWR VGND sg13g2_nand2_1
X_3298_ net992 net1062 _1736_ VPWR VGND sg13g2_nor2b_1
XFILLER_38_461 VPWR VGND sg13g2_decap_8
XFILLER_26_656 VPWR VGND sg13g2_fill_1
XFILLER_40_114 VPWR VGND sg13g2_decap_8
XFILLER_15_56 VPWR VGND sg13g2_decap_4
X_5939_ s0.data_out\[8\]\[7\] s0.data_out\[7\]\[7\] net1021 _1553_ VPWR VGND sg13g2_mux2_1
XFILLER_15_67 VPWR VGND sg13g2_fill_1
XFILLER_40_169 VPWR VGND sg13g2_fill_2
X_6104__173 VPWR VGND net173 sg13g2_tiehi
XFILLER_1_711 VPWR VGND sg13g2_decap_8
Xoutput9 net9 uo_out[7] VPWR VGND sg13g2_buf_1
XFILLER_49_737 VPWR VGND sg13g2_decap_8
XFILLER_1_788 VPWR VGND sg13g2_decap_8
XFILLER_45_921 VPWR VGND sg13g2_decap_8
X_6111__166 VPWR VGND net166 sg13g2_tiehi
XFILLER_45_998 VPWR VGND sg13g2_decap_8
XFILLER_44_453 VPWR VGND sg13g2_fill_2
XFILLER_44_442 VPWR VGND sg13g2_decap_8
XFILLER_17_678 VPWR VGND sg13g2_fill_2
XFILLER_16_177 VPWR VGND sg13g2_fill_1
XFILLER_9_800 VPWR VGND sg13g2_decap_8
XFILLER_9_811 VPWR VGND sg13g2_fill_1
XFILLER_9_844 VPWR VGND sg13g2_fill_2
XFILLER_4_560 VPWR VGND sg13g2_fill_2
X_4270_ _2610_ net1246 _2609_ VPWR VGND sg13g2_nand2_1
X_3221_ _1665_ net1002 _1617_ _1666_ VPWR VGND sg13g2_a21o_1
XFILLER_39_214 VPWR VGND sg13g2_fill_2
X_3152_ net1002 net1071 _1604_ VPWR VGND sg13g2_nor2b_1
XFILLER_39_269 VPWR VGND sg13g2_fill_2
XFILLER_27_409 VPWR VGND sg13g2_decap_8
XFILLER_47_280 VPWR VGND sg13g2_fill_2
XFILLER_36_987 VPWR VGND sg13g2_decap_8
XFILLER_22_136 VPWR VGND sg13g2_decap_8
X_3985_ net1281 _2357_ _2358_ VPWR VGND sg13g2_nor2b_1
X_5724_ s0.data_out\[8\]\[0\] s0.data_out\[9\]\[0\] net1041 _1358_ VPWR VGND sg13g2_mux2_1
X_5655_ VGND VPWR net1036 _1299_ _1300_ _1249_ sg13g2_a21oi_1
X_4606_ VGND VPWR net1158 s0.data_out\[17\]\[6\] _0349_ _0348_ sg13g2_a21oi_1
XFILLER_11_1023 VPWR VGND sg13g2_decap_4
Xhold310 s0.data_new_delayed\[0\] VPWR VGND net606 sg13g2_dlygate4sd3_1
X_5586_ s0.data_out\[9\]\[0\] s0.data_out\[10\]\[0\] net1084 _1239_ VPWR VGND sg13g2_mux2_1
X_4537_ _0290_ _0289_ _0273_ VPWR VGND sg13g2_nand2b_1
X_6058__223 VPWR VGND net223 sg13g2_tiehi
X_4468_ net1289 VPWR _2787_ VGND net927 _2786_ sg13g2_o21ai_1
X_6207_ net273 VGND VPWR _0257_ s0.data_out\[1\]\[7\] clknet_leaf_10_clk sg13g2_dfrbpq_2
X_3419_ VGND VPWR _1846_ net581 net1311 sg13g2_or2_1
X_6138_ net137 VGND VPWR net466 s0.was_valid_out\[6\][0] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_4399_ _2727_ net1196 _2726_ VPWR VGND sg13g2_nand2b_1
XFILLER_39_770 VPWR VGND sg13g2_decap_4
X_6069_ net211 VGND VPWR _0119_ s0.shift_out\[12\][0] clknet_leaf_27_clk sg13g2_dfrbpq_1
XFILLER_18_409 VPWR VGND sg13g2_fill_2
XFILLER_26_22 VPWR VGND sg13g2_decap_8
XFILLER_42_957 VPWR VGND sg13g2_decap_8
X_5991__23 VPWR VGND net23 sg13g2_tiehi
XFILLER_13_125 VPWR VGND sg13g2_fill_2
XFILLER_6_869 VPWR VGND sg13g2_fill_2
XFILLER_3_59 VPWR VGND sg13g2_fill_2
XFILLER_3_48 VPWR VGND sg13g2_decap_8
XFILLER_1_585 VPWR VGND sg13g2_decap_8
XFILLER_49_534 VPWR VGND sg13g2_decap_8
XFILLER_37_718 VPWR VGND sg13g2_decap_8
XFILLER_18_987 VPWR VGND sg13g2_decap_8
XFILLER_45_795 VPWR VGND sg13g2_decap_8
XFILLER_32_412 VPWR VGND sg13g2_decap_8
X_3770_ net1298 net300 _0235_ VPWR VGND sg13g2_and2_1
XFILLER_34_1012 VPWR VGND sg13g2_decap_8
XFILLER_13_681 VPWR VGND sg13g2_fill_2
XFILLER_13_692 VPWR VGND sg13g2_fill_2
X_5440_ _1082_ _1094_ _1107_ _1108_ _1109_ VPWR VGND sg13g2_or4_1
X_5371_ net1092 net1055 _1043_ VPWR VGND sg13g2_nor2b_1
X_4322_ VGND VPWR _2584_ _2654_ _2655_ net1193 sg13g2_a21oi_1
X_4253_ _2592_ net1192 _2564_ _2593_ VPWR VGND sg13g2_a21o_1
X_3204_ VPWR _0185_ net518 VGND sg13g2_inv_1
X_4184_ net1202 VPWR _2530_ VGND _2528_ _2529_ sg13g2_o21ai_1
X_3135_ _1590_ _1587_ _1589_ VPWR VGND sg13g2_nand2_1
XFILLER_28_718 VPWR VGND sg13g2_fill_2
XFILLER_24_979 VPWR VGND sg13g2_decap_8
X_3968_ net944 net1045 _2342_ VPWR VGND sg13g2_nor2b_1
X_5707_ VGND VPWR net1223 net1214 _0148_ _1346_ sg13g2_a21oi_1
X_3899_ net1291 net306 _0247_ VPWR VGND sg13g2_and2_1
X_5638_ net1346 VPWR _1285_ VGND net934 _1284_ sg13g2_o21ai_1
XFILLER_12_68 VPWR VGND sg13g2_decap_8
XFILLER_3_817 VPWR VGND sg13g2_decap_8
X_5569_ _1207_ _1209_ _1226_ VPWR VGND sg13g2_nor2b_1
XFILLER_2_327 VPWR VGND sg13g2_decap_8
Xhold162 s0.data_out\[1\]\[2\] VPWR VGND net458 sg13g2_dlygate4sd3_1
Xhold151 _2203_ VPWR VGND net447 sg13g2_dlygate4sd3_1
Xhold140 s0.data_out\[10\]\[3\] VPWR VGND net436 sg13g2_dlygate4sd3_1
Xhold195 s0.data_out\[2\]\[6\] VPWR VGND net491 sg13g2_dlygate4sd3_1
Xhold184 s0.data_out\[17\]\[3\] VPWR VGND net480 sg13g2_dlygate4sd3_1
Xhold173 s0.data_out\[20\]\[4\] VPWR VGND net469 sg13g2_dlygate4sd3_1
XFILLER_37_32 VPWR VGND sg13g2_decap_4
XFILLER_33_209 VPWR VGND sg13g2_decap_4
XFILLER_27_784 VPWR VGND sg13g2_decap_4
XFILLER_42_743 VPWR VGND sg13g2_decap_4
XFILLER_6_677 VPWR VGND sg13g2_fill_1
XFILLER_6_666 VPWR VGND sg13g2_decap_8
XFILLER_5_154 VPWR VGND sg13g2_decap_8
XFILLER_5_132 VPWR VGND sg13g2_fill_2
XFILLER_2_861 VPWR VGND sg13g2_decap_8
XFILLER_38_7 VPWR VGND sg13g2_fill_2
XFILLER_37_537 VPWR VGND sg13g2_fill_1
XFILLER_18_740 VPWR VGND sg13g2_fill_1
X_4940_ net1122 s0.data_out\[14\]\[0\] _0653_ VPWR VGND sg13g2_and2_1
X_4871_ VGND VPWR _0589_ net591 net1318 sg13g2_or2_1
X_6048__233 VPWR VGND net233 sg13g2_tiehi
XFILLER_17_294 VPWR VGND sg13g2_fill_1
X_3822_ VPWR _0242_ _2210_ VGND sg13g2_inv_1
XFILLER_21_927 VPWR VGND sg13g2_decap_8
X_3753_ _2150_ net971 _2149_ VPWR VGND sg13g2_nand2b_1
X_3684_ net1307 VPWR _2086_ VGND net932 _2085_ sg13g2_o21ai_1
X_5423_ VGND VPWR _1092_ _1086_ net1236 sg13g2_or2_1
X_5354_ _1028_ net938 _1027_ VPWR VGND sg13g2_nand2_1
X_4305_ s0.data_out\[19\]\[1\] s0.data_out\[20\]\[1\] net1199 _2640_ VPWR VGND sg13g2_mux2_1
X_6055__226 VPWR VGND net226 sg13g2_tiehi
X_5285_ s0.data_out\[13\]\[7\] s0.data_out\[12\]\[7\] net1111 _0966_ VPWR VGND sg13g2_mux2_1
X_4236_ _2576_ net1203 _2575_ VPWR VGND sg13g2_nand2b_1
X_4167_ net1190 s0.data_out\[20\]\[0\] _2515_ VPWR VGND sg13g2_and2_1
X_3118_ net1252 _1572_ _1575_ VPWR VGND sg13g2_nor2_1
X_4098_ VPWR _2457_ net1203 VGND sg13g2_inv_1
XFILLER_36_581 VPWR VGND sg13g2_decap_4
XFILLER_23_67 VPWR VGND sg13g2_fill_2
XFILLER_3_4 VPWR VGND sg13g2_fill_2
XFILLER_24_1000 VPWR VGND sg13g2_decap_8
XFILLER_47_857 VPWR VGND sg13g2_decap_8
XFILLER_19_548 VPWR VGND sg13g2_fill_1
XFILLER_46_367 VPWR VGND sg13g2_decap_8
XFILLER_46_378 VPWR VGND sg13g2_fill_1
XFILLER_27_570 VPWR VGND sg13g2_fill_1
XFILLER_14_231 VPWR VGND sg13g2_fill_2
XFILLER_27_592 VPWR VGND sg13g2_decap_8
XFILLER_42_573 VPWR VGND sg13g2_fill_1
XFILLER_42_562 VPWR VGND sg13g2_decap_8
XFILLER_11_960 VPWR VGND sg13g2_decap_8
XFILLER_30_768 VPWR VGND sg13g2_decap_8
XFILLER_7_964 VPWR VGND sg13g2_decap_8
XFILLER_9_1027 VPWR VGND sg13g2_fill_2
X_5070_ s0.data_out\[13\]\[0\] s0.data_out\[14\]\[0\] net1131 _0771_ VPWR VGND sg13g2_mux2_1
X_4021_ _2388_ VPWR _2394_ VGND _2383_ _2390_ sg13g2_o21ai_1
X_5972_ net44 VGND VPWR _0022_ s0.data_out\[20\]\[7\] clknet_leaf_0_clk sg13g2_dfrbpq_2
X_4923_ VGND VPWR _0640_ net1209 net310 sg13g2_or2_1
XFILLER_33_551 VPWR VGND sg13g2_fill_1
X_4854_ net1149 VPWR _0574_ VGND _0572_ _0573_ sg13g2_o21ai_1
X_4785_ VGND VPWR net1161 _0513_ _0514_ _0457_ sg13g2_a21oi_1
XFILLER_20_256 VPWR VGND sg13g2_fill_2
X_3805_ _2195_ VPWR _2196_ VGND _2191_ _2194_ sg13g2_o21ai_1
X_3736_ VGND VPWR net971 _2132_ _2133_ _2083_ sg13g2_a21oi_1
X_3667_ net959 net1072 _2071_ VPWR VGND sg13g2_nor2b_1
XFILLER_47_1011 VPWR VGND sg13g2_decap_8
X_5406_ VPWR VGND _1007_ net1282 _1073_ net1279 _1075_ _1070_ sg13g2_a221oi_1
X_3598_ _1952_ _2006_ _2007_ VPWR VGND sg13g2_and2_1
XFILLER_0_628 VPWR VGND sg13g2_decap_8
X_5337_ _1013_ s0.data_out\[11\]\[1\] net1109 VPWR VGND sg13g2_nand2b_1
X_5268_ s0.data_out\[13\]\[1\] s0.data_out\[12\]\[1\] net1108 _0949_ VPWR VGND sg13g2_mux2_1
X_4219_ net1204 _2559_ _2560_ _2561_ VPWR VGND sg13g2_nor3_1
X_5199_ s0.data_out\[12\]\[0\] s0.data_out\[13\]\[0\] net1120 _0888_ VPWR VGND sg13g2_mux2_1
XFILLER_18_12 VPWR VGND sg13g2_decap_8
XFILLER_37_890 VPWR VGND sg13g2_fill_2
XFILLER_11_245 VPWR VGND sg13g2_decap_8
XFILLER_4_956 VPWR VGND sg13g2_decap_8
Xfanout1212 _2480_ net1212 VPWR VGND sg13g2_buf_8
Xfanout1201 s0.valid_out\[20\][0] net1201 VPWR VGND sg13g2_buf_2
Xfanout1223 uio_in[1] net1223 VPWR VGND sg13g2_buf_8
Xfanout1245 ui_in[6] net1245 VPWR VGND sg13g2_buf_8
Xfanout1256 net1259 net1256 VPWR VGND sg13g2_buf_8
Xfanout1234 ui_in[7] net1234 VPWR VGND sg13g2_buf_8
Xfanout1289 net1290 net1289 VPWR VGND sg13g2_buf_8
XFILLER_19_301 VPWR VGND sg13g2_fill_2
Xfanout1278 net1279 net1278 VPWR VGND sg13g2_buf_8
Xfanout1267 ui_in[3] net1267 VPWR VGND sg13g2_buf_8
XFILLER_47_654 VPWR VGND sg13g2_decap_8
XFILLER_46_175 VPWR VGND sg13g2_decap_4
XFILLER_35_849 VPWR VGND sg13g2_fill_2
XFILLER_35_816 VPWR VGND sg13g2_decap_8
XFILLER_19_378 VPWR VGND sg13g2_decap_4
XFILLER_19_389 VPWR VGND sg13g2_fill_1
XFILLER_34_315 VPWR VGND sg13g2_fill_2
X_4570_ VPWR _0040_ net494 VGND sg13g2_inv_1
X_3521_ net972 _1934_ _1940_ VPWR VGND sg13g2_nor2_1
XFILLER_6_260 VPWR VGND sg13g2_fill_1
X_3452_ _1874_ VPWR _1875_ VGND _1870_ _1873_ sg13g2_o21ai_1
X_6171_ net101 VGND VPWR _0221_ s0.data_out\[4\]\[7\] clknet_leaf_12_clk sg13g2_dfrbpq_2
XFILLER_41_2 VPWR VGND sg13g2_fill_1
X_3383_ VGND VPWR _1816_ net1209 net309 sg13g2_or2_1
X_5122_ net1333 VPWR _0817_ VGND net937 _0816_ sg13g2_o21ai_1
X_6052__229 VPWR VGND net229 sg13g2_tiehi
XFILLER_27_0 VPWR VGND sg13g2_decap_4
XFILLER_38_621 VPWR VGND sg13g2_fill_1
X_5053_ _0740_ _0757_ _0758_ VPWR VGND sg13g2_nor2b_1
X_4004_ VGND VPWR _2377_ _2371_ net1232 sg13g2_or2_1
XFILLER_38_676 VPWR VGND sg13g2_fill_1
XFILLER_37_164 VPWR VGND sg13g2_fill_2
XFILLER_26_827 VPWR VGND sg13g2_fill_1
X_5955_ net62 VGND VPWR _0005_ s0.data_out\[21\]\[2\] clknet_leaf_37_clk sg13g2_dfrbpq_1
XFILLER_40_318 VPWR VGND sg13g2_fill_2
X_4906_ VGND VPWR net1137 _0622_ _0623_ _0573_ sg13g2_a21oi_1
X_5886_ VPWR _0169_ _1504_ VGND sg13g2_inv_1
X_4837_ VGND VPWR net1134 net387 _0559_ _0558_ sg13g2_a21oi_1
XFILLER_14_1010 VPWR VGND sg13g2_decap_8
X_4768_ s0.data_out\[17\]\[6\] s0.data_out\[16\]\[6\] net1154 _0497_ VPWR VGND sg13g2_mux2_1
X_3719_ VPWR _0233_ net516 VGND sg13g2_inv_1
X_4699_ VPWR _0052_ net497 VGND sg13g2_inv_1
XFILLER_49_919 VPWR VGND sg13g2_decap_8
Xhold22 s0.genblk1\[5\].modules.bubble VPWR VGND net318 sg13g2_dlygate4sd3_1
Xhold11 s0.genblk1\[8\].modules.bubble VPWR VGND net307 sg13g2_dlygate4sd3_1
XFILLER_48_429 VPWR VGND sg13g2_decap_8
Xhold33 _0248_ VPWR VGND net329 sg13g2_dlygate4sd3_1
Xhold44 net1014 VPWR VGND net340 sg13g2_dlygate4sd3_1
Xhold55 s0.data_out\[0\]\[6\] VPWR VGND net351 sg13g2_dlygate4sd3_1
Xhold88 _0200_ VPWR VGND net384 sg13g2_dlygate4sd3_1
Xhold77 _0001_ VPWR VGND net373 sg13g2_dlygate4sd3_1
Xhold99 s0.data_out\[20\]\[5\] VPWR VGND net395 sg13g2_dlygate4sd3_1
XFILLER_21_1025 VPWR VGND sg13g2_decap_4
Xhold66 _0008_ VPWR VGND net362 sg13g2_dlygate4sd3_1
XFILLER_29_88 VPWR VGND sg13g2_fill_1
XFILLER_28_131 VPWR VGND sg13g2_fill_2
XFILLER_45_32 VPWR VGND sg13g2_fill_1
XFILLER_25_860 VPWR VGND sg13g2_decap_4
XFILLER_43_178 VPWR VGND sg13g2_decap_8
XFILLER_40_852 VPWR VGND sg13g2_decap_4
XFILLER_12_554 VPWR VGND sg13g2_decap_4
XFILLER_40_874 VPWR VGND sg13g2_fill_2
XFILLER_4_753 VPWR VGND sg13g2_fill_1
XFILLER_4_742 VPWR VGND sg13g2_decap_8
XFILLER_4_775 VPWR VGND sg13g2_decap_4
Xfanout1020 net1021 net1020 VPWR VGND sg13g2_buf_8
Xfanout1031 net1034 net1031 VPWR VGND sg13g2_buf_8
Xfanout1042 net1044 net1042 VPWR VGND sg13g2_buf_1
XFILLER_0_992 VPWR VGND sg13g2_decap_8
Xfanout1053 net1056 net1053 VPWR VGND sg13g2_buf_8
Xfanout1064 net604 net1064 VPWR VGND sg13g2_buf_8
XFILLER_48_941 VPWR VGND sg13g2_decap_8
Xfanout1086 net1087 net1086 VPWR VGND sg13g2_buf_1
Xfanout1075 net1076 net1075 VPWR VGND sg13g2_buf_2
Xfanout1097 net1098 net1097 VPWR VGND sg13g2_buf_8
XFILLER_35_602 VPWR VGND sg13g2_fill_2
XFILLER_35_646 VPWR VGND sg13g2_fill_1
XFILLER_19_197 VPWR VGND sg13g2_fill_1
X_5740_ s0.data_out\[8\]\[2\] s0.data_out\[9\]\[2\] net1041 _1372_ VPWR VGND sg13g2_mux2_1
X_5671_ _1315_ net1039 _1290_ _1316_ VPWR VGND sg13g2_a21o_1
X_4622_ VGND VPWR net1169 _0362_ _0363_ _0319_ sg13g2_a21oi_1
X_4553_ _0302_ _0303_ _0037_ VPWR VGND sg13g2_nor2_1
X_4484_ net1288 VPWR _2801_ VGND net926 _2800_ sg13g2_o21ai_1
X_3504_ _1856_ _1917_ net1258 _1925_ VPWR VGND sg13g2_nand3_1
X_3435_ _1856_ _1859_ net1312 _1860_ VPWR VGND sg13g2_nand3_1
XFILLER_44_1025 VPWR VGND sg13g2_decap_4
X_3366_ s0.data_out\[6\]\[5\] s0.data_out\[5\]\[5\] net998 _1799_ VPWR VGND sg13g2_mux2_1
X_6154_ net119 VGND VPWR _0204_ s0.data_out\[5\]\[2\] clknet_leaf_5_clk sg13g2_dfrbpq_2
X_5105_ VGND VPWR net1115 net430 _0802_ _0801_ sg13g2_a21oi_1
X_6085_ net193 VGND VPWR _0135_ s0.data_out\[10\]\[0\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_3297_ net992 s0.data_out\[5\]\[3\] _1735_ VPWR VGND sg13g2_and2_1
X_5036_ VPWR _0741_ _0740_ VGND sg13g2_inv_1
XFILLER_13_307 VPWR VGND sg13g2_fill_2
XFILLER_41_627 VPWR VGND sg13g2_decap_4
X_5938_ _1552_ net1020 net517 VPWR VGND sg13g2_nand2_1
XFILLER_13_329 VPWR VGND sg13g2_decap_8
X_5869_ _1489_ VPWR _1490_ VGND _1485_ _1488_ sg13g2_o21ai_1
XFILLER_49_716 VPWR VGND sg13g2_decap_8
XFILLER_0_222 VPWR VGND sg13g2_decap_8
XFILLER_1_767 VPWR VGND sg13g2_decap_8
XFILLER_45_900 VPWR VGND sg13g2_decap_8
XFILLER_29_451 VPWR VGND sg13g2_fill_1
XFILLER_45_977 VPWR VGND sg13g2_decap_8
XFILLER_32_605 VPWR VGND sg13g2_fill_1
XFILLER_31_137 VPWR VGND sg13g2_decap_4
XFILLER_40_660 VPWR VGND sg13g2_decap_4
XFILLER_8_300 VPWR VGND sg13g2_decap_4
XFILLER_9_823 VPWR VGND sg13g2_fill_1
XFILLER_40_693 VPWR VGND sg13g2_fill_2
XFILLER_12_395 VPWR VGND sg13g2_fill_1
X_3220_ s0.data_out\[7\]\[3\] s0.data_out\[6\]\[3\] net1011 _1665_ VPWR VGND sg13g2_mux2_1
X_3151_ net1001 s0.data_out\[6\]\[1\] _1603_ VPWR VGND sg13g2_and2_1
XFILLER_35_432 VPWR VGND sg13g2_decap_4
XFILLER_36_966 VPWR VGND sg13g2_decap_8
X_3984_ _2292_ VPWR _2357_ VGND net928 _2356_ sg13g2_o21ai_1
X_5723_ net1221 _1352_ _0153_ VPWR VGND sg13g2_nor2_1
XFILLER_31_671 VPWR VGND sg13g2_fill_1
X_5654_ s0.data_out\[10\]\[1\] s0.data_out\[9\]\[1\] net1041 _1299_ VPWR VGND sg13g2_mux2_1
XFILLER_11_1002 VPWR VGND sg13g2_decap_8
X_4605_ net1158 net1050 _0348_ VPWR VGND sg13g2_nor2b_1
Xhold300 _1532_ VPWR VGND net596 sg13g2_dlygate4sd3_1
Xhold311 s0.data_new_delayed\[5\] VPWR VGND net607 sg13g2_dlygate4sd3_1
X_5585_ net1221 _1233_ _0134_ VPWR VGND sg13g2_nor2_1
X_4536_ _0278_ VPWR _0289_ VGND _0282_ _0284_ sg13g2_o21ai_1
X_4467_ VGND VPWR net1172 net570 _2786_ _2785_ sg13g2_a21oi_1
X_5997__289 VPWR VGND net289 sg13g2_tiehi
X_6206_ net286 VGND VPWR _0256_ s0.data_out\[1\]\[6\] clknet_leaf_10_clk sg13g2_dfrbpq_2
X_4398_ VGND VPWR net1183 _2725_ _2726_ _2671_ sg13g2_a21oi_1
X_3418_ net1311 VPWR _1845_ VGND net915 _1844_ sg13g2_o21ai_1
X_6137_ net138 VGND VPWR _0187_ s0.genblk1\[6\].modules.bubble clknet_leaf_13_clk
+ sg13g2_dfrbpq_1
X_3349_ VGND VPWR net992 _1781_ _1782_ _1736_ sg13g2_a21oi_1
XFILLER_46_719 VPWR VGND sg13g2_decap_8
X_6068_ net212 VGND VPWR _0118_ s0.data_out\[12\]\[7\] clknet_leaf_26_clk sg13g2_dfrbpq_2
XFILLER_38_270 VPWR VGND sg13g2_decap_4
X_5019_ VGND VPWR net1124 _0723_ _0724_ _0674_ sg13g2_a21oi_1
XFILLER_26_56 VPWR VGND sg13g2_decap_4
XFILLER_27_988 VPWR VGND sg13g2_decap_8
XFILLER_42_936 VPWR VGND sg13g2_decap_8
XFILLER_14_627 VPWR VGND sg13g2_decap_4
XFILLER_41_446 VPWR VGND sg13g2_decap_8
XFILLER_10_800 VPWR VGND sg13g2_fill_1
XFILLER_42_55 VPWR VGND sg13g2_decap_4
XFILLER_10_866 VPWR VGND sg13g2_fill_2
XFILLER_21_192 VPWR VGND sg13g2_decap_4
XFILLER_5_347 VPWR VGND sg13g2_fill_1
XFILLER_5_336 VPWR VGND sg13g2_decap_8
XFILLER_49_513 VPWR VGND sg13g2_decap_8
XFILLER_1_564 VPWR VGND sg13g2_decap_8
XFILLER_29_270 VPWR VGND sg13g2_fill_2
XFILLER_18_966 VPWR VGND sg13g2_decap_8
XFILLER_29_292 VPWR VGND sg13g2_fill_2
XFILLER_45_774 VPWR VGND sg13g2_decap_8
XFILLER_44_284 VPWR VGND sg13g2_fill_2
XFILLER_33_969 VPWR VGND sg13g2_decap_8
XFILLER_20_608 VPWR VGND sg13g2_decap_8
XFILLER_8_163 VPWR VGND sg13g2_decap_4
XFILLER_9_675 VPWR VGND sg13g2_fill_2
X_5370_ VGND VPWR _0983_ _1041_ _1042_ net1105 sg13g2_a21oi_1
X_4321_ _2654_ s0.data_out\[19\]\[3\] net1199 VPWR VGND sg13g2_nand2b_1
XFILLER_5_881 VPWR VGND sg13g2_decap_8
X_4252_ s0.data_out\[21\]\[7\] s0.data_out\[20\]\[7\] net1198 _2592_ VPWR VGND sg13g2_mux2_1
X_3203_ _1648_ VPWR _1649_ VGND _1644_ _1647_ sg13g2_o21ai_1
XFILLER_41_1028 VPWR VGND sg13g2_fill_1
XFILLER_41_1017 VPWR VGND sg13g2_decap_8
X_4183_ net1191 net1065 _2529_ VPWR VGND sg13g2_nor2b_1
X_3134_ _2468_ VPWR _1589_ VGND s0.was_valid_out\[6\][0] net1020 sg13g2_o21ai_1
XFILLER_24_903 VPWR VGND sg13g2_fill_1
XFILLER_36_785 VPWR VGND sg13g2_decap_4
XFILLER_35_251 VPWR VGND sg13g2_decap_8
X_3967_ VGND VPWR _2252_ _2340_ _2341_ net952 sg13g2_a21oi_1
XFILLER_10_129 VPWR VGND sg13g2_decap_8
X_5706_ net1224 net1057 _1346_ VPWR VGND sg13g2_nor2_1
X_3898_ VGND VPWR _2277_ _2281_ _0246_ _2282_ sg13g2_a21oi_1
Xclkbuf_leaf_30_clk clknet_3_4__leaf_clk clknet_leaf_30_clk VPWR VGND sg13g2_buf_8
XFILLER_31_490 VPWR VGND sg13g2_fill_2
X_5637_ VGND VPWR net1038 s0.data_out\[9\]\[6\] _1284_ _1283_ sg13g2_a21oi_1
X_5568_ _1210_ _1218_ _1220_ _1225_ VPWR VGND sg13g2_nor3_1
X_4519_ VGND VPWR _0272_ _2828_ net1231 sg13g2_or2_1
X_6101__177 VPWR VGND net177 sg13g2_tiehi
Xhold141 s0.data_out\[3\]\[0\] VPWR VGND net437 sg13g2_dlygate4sd3_1
Xhold152 s0.data_out\[1\]\[0\] VPWR VGND net448 sg13g2_dlygate4sd3_1
Xhold130 s0.data_out\[2\]\[1\] VPWR VGND net426 sg13g2_dlygate4sd3_1
Xhold174 s0.data_out\[4\]\[5\] VPWR VGND net470 sg13g2_dlygate4sd3_1
Xhold185 s0.data_out\[10\]\[5\] VPWR VGND net481 sg13g2_dlygate4sd3_1
X_5499_ VPWR _0127_ _1159_ VGND sg13g2_inv_1
Xhold163 _2311_ VPWR VGND net459 sg13g2_dlygate4sd3_1
Xhold196 _2224_ VPWR VGND net492 sg13g2_dlygate4sd3_1
XFILLER_46_527 VPWR VGND sg13g2_decap_8
XFILLER_37_55 VPWR VGND sg13g2_decap_8
XFILLER_2_1022 VPWR VGND sg13g2_decap_8
XFILLER_15_903 VPWR VGND sg13g2_fill_2
XFILLER_26_240 VPWR VGND sg13g2_decap_8
XFILLER_14_413 VPWR VGND sg13g2_fill_2
XFILLER_15_936 VPWR VGND sg13g2_fill_2
XFILLER_27_774 VPWR VGND sg13g2_decap_4
XFILLER_18_1008 VPWR VGND sg13g2_decap_8
XFILLER_14_479 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_21_clk clknet_3_7__leaf_clk clknet_leaf_21_clk VPWR VGND sg13g2_buf_8
XFILLER_2_840 VPWR VGND sg13g2_decap_8
XFILLER_49_332 VPWR VGND sg13g2_decap_4
XFILLER_49_387 VPWR VGND sg13g2_decap_8
XFILLER_18_763 VPWR VGND sg13g2_fill_1
XFILLER_17_240 VPWR VGND sg13g2_fill_1
X_4870_ net1317 VPWR _0588_ VGND net922 _0587_ sg13g2_o21ai_1
X_3821_ _2209_ VPWR _2210_ VGND net1298 net417 sg13g2_o21ai_1
Xclkbuf_leaf_12_clk clknet_3_3__leaf_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
X_3752_ VGND VPWR net960 _2148_ _2149_ _2092_ sg13g2_a21oi_1
XFILLER_9_494 VPWR VGND sg13g2_fill_2
X_3683_ VGND VPWR net960 net446 _2085_ _2084_ sg13g2_a21oi_1
X_5422_ _1091_ _1090_ net1242 _1086_ net1236 VPWR VGND sg13g2_a22oi_1
X_5353_ s0.data_out\[11\]\[3\] s0.data_out\[12\]\[3\] net1108 _1027_ VPWR VGND sg13g2_mux2_1
X_4304_ VPWR _0015_ _2639_ VGND sg13g2_inv_1
X_5284_ _0965_ net1110 net594 VPWR VGND sg13g2_nand2_1
X_4235_ VGND VPWR net1190 _2574_ _2575_ _2522_ sg13g2_a21oi_1
X_4166_ net1190 net1073 _2514_ VPWR VGND sg13g2_nor2b_1
X_3117_ _1567_ _1506_ net1256 _1574_ VPWR VGND sg13g2_a21o_1
X_4097_ _2456_ net1194 VPWR VGND sg13g2_inv_2
XFILLER_24_711 VPWR VGND sg13g2_fill_2
XFILLER_23_210 VPWR VGND sg13g2_decap_8
XFILLER_24_766 VPWR VGND sg13g2_decap_8
XFILLER_24_777 VPWR VGND sg13g2_fill_2
X_4999_ VGND VPWR _0705_ net554 net1318 sg13g2_or2_1
XFILLER_23_276 VPWR VGND sg13g2_fill_2
XFILLER_7_409 VPWR VGND sg13g2_fill_1
XFILLER_11_449 VPWR VGND sg13g2_fill_2
XFILLER_20_983 VPWR VGND sg13g2_decap_8
XFILLER_48_21 VPWR VGND sg13g2_decap_8
XFILLER_47_836 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_fill_2
XFILLER_34_508 VPWR VGND sg13g2_decap_4
XFILLER_15_722 VPWR VGND sg13g2_fill_2
XFILLER_9_15 VPWR VGND sg13g2_fill_2
XFILLER_9_59 VPWR VGND sg13g2_decap_8
XFILLER_7_943 VPWR VGND sg13g2_decap_8
XFILLER_31_1027 VPWR VGND sg13g2_fill_2
XFILLER_6_464 VPWR VGND sg13g2_fill_2
XFILLER_9_1006 VPWR VGND sg13g2_decap_8
XFILLER_38_803 VPWR VGND sg13g2_fill_2
X_4020_ _2379_ _2389_ _2391_ _2392_ _2393_ VPWR VGND sg13g2_and4_1
Xclkbuf_leaf_1_clk clknet_3_0__leaf_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
XFILLER_38_825 VPWR VGND sg13g2_decap_8
XFILLER_37_357 VPWR VGND sg13g2_decap_8
XFILLER_46_880 VPWR VGND sg13g2_decap_8
X_5971_ net45 VGND VPWR _0021_ s0.data_out\[20\]\[6\] clknet_leaf_0_clk sg13g2_dfrbpq_2
X_4922_ _0527_ _0528_ _0637_ _0638_ _0639_ VPWR VGND sg13g2_nor4_1
X_4853_ net1136 net1055 _0573_ VPWR VGND sg13g2_nor2b_1
X_4784_ _0512_ net1147 _0458_ _0513_ VPWR VGND sg13g2_a21o_1
XFILLER_20_235 VPWR VGND sg13g2_decap_8
X_3804_ VGND VPWR _2195_ net488 net1297 sg13g2_or2_1
X_3735_ _2131_ net960 _2084_ _2132_ VPWR VGND sg13g2_a21o_1
X_5405_ net1279 _1070_ _1074_ VPWR VGND sg13g2_nor2_1
X_3666_ net960 s0.data_out\[2\]\[1\] _2070_ VPWR VGND sg13g2_and2_1
X_3597_ _2006_ net980 _2005_ VPWR VGND sg13g2_nand2b_1
XFILLER_0_607 VPWR VGND sg13g2_decap_8
X_5336_ VPWR _0111_ _1012_ VGND sg13g2_inv_1
X_5267_ _0948_ net1109 net528 VPWR VGND sg13g2_nand2_1
X_4218_ s0.valid_out\[21\][0] s0.data_out\[20\]\[6\] _2560_ VPWR VGND sg13g2_nor2_1
X_5198_ net1220 _0880_ _0881_ _0098_ VPWR VGND sg13g2_nor3_1
XFILLER_29_836 VPWR VGND sg13g2_decap_8
XFILLER_18_68 VPWR VGND sg13g2_fill_2
X_4149_ VGND VPWR _2474_ net912 net8 _2501_ sg13g2_a21oi_1
XFILLER_28_346 VPWR VGND sg13g2_decap_8
XFILLER_28_357 VPWR VGND sg13g2_fill_2
XFILLER_29_869 VPWR VGND sg13g2_fill_2
XFILLER_24_541 VPWR VGND sg13g2_decap_8
Xclkload0 clknet_3_3__leaf_clk clkload0/X VPWR VGND sg13g2_buf_8
XFILLER_4_935 VPWR VGND sg13g2_decap_8
Xfanout1213 _2480_ net1213 VPWR VGND sg13g2_buf_8
Xfanout1202 net1203 net1202 VPWR VGND sg13g2_buf_8
X_6038__244 VPWR VGND net244 sg13g2_tiehi
Xfanout1246 net1249 net1246 VPWR VGND sg13g2_buf_8
Xfanout1224 uio_in[1] net1224 VPWR VGND sg13g2_buf_1
Xfanout1235 net1238 net1235 VPWR VGND sg13g2_buf_8
Xfanout1257 net1259 net1257 VPWR VGND sg13g2_buf_1
Xfanout1268 net1272 net1268 VPWR VGND sg13g2_buf_8
Xfanout1279 net1280 net1279 VPWR VGND sg13g2_buf_8
XFILLER_47_633 VPWR VGND sg13g2_decap_8
X_6045__237 VPWR VGND net237 sg13g2_tiehi
XFILLER_15_596 VPWR VGND sg13g2_fill_1
X_3520_ net319 net978 _1939_ VPWR VGND sg13g2_nor2_1
X_3451_ VGND VPWR _1874_ net538 net1313 sg13g2_or2_1
X_6170_ net102 VGND VPWR _0220_ s0.data_out\[4\]\[6\] clknet_leaf_12_clk sg13g2_dfrbpq_2
X_3382_ _1706_ _1813_ _1814_ _1815_ VPWR VGND sg13g2_nor3_1
X_5121_ VGND VPWR net1114 net597 _0816_ _0815_ sg13g2_a21oi_1
X_5052_ _0751_ VPWR _0757_ VGND _0746_ _0753_ sg13g2_o21ai_1
X_4003_ VGND VPWR _2376_ _2374_ net1241 sg13g2_or2_1
XFILLER_1_82 VPWR VGND sg13g2_decap_4
Xheichips25_top_sorter_20 VPWR VGND uio_out[5] sg13g2_tielo
XFILLER_25_316 VPWR VGND sg13g2_fill_2
XFILLER_37_198 VPWR VGND sg13g2_decap_4
X_5954_ net63 VGND VPWR _0004_ s0.data_out\[21\]\[1\] clknet_leaf_37_clk sg13g2_dfrbpq_1
X_4905_ s0.data_out\[16\]\[5\] s0.data_out\[15\]\[5\] net1143 _0622_ VPWR VGND sg13g2_mux2_1
XFILLER_33_360 VPWR VGND sg13g2_fill_2
X_5885_ _1503_ VPWR _1504_ VGND net1327 net434 sg13g2_o21ai_1
XFILLER_34_894 VPWR VGND sg13g2_decap_8
X_4836_ net1134 net1062 _0558_ VPWR VGND sg13g2_nor2b_1
XFILLER_21_533 VPWR VGND sg13g2_fill_2
X_4767_ _0496_ net1152 net546 VPWR VGND sg13g2_nand2_1
X_3718_ _2115_ VPWR _2116_ VGND _2111_ _2114_ sg13g2_o21ai_1
X_4698_ _0433_ VPWR _0434_ VGND _0429_ _0432_ sg13g2_o21ai_1
XFILLER_20_14 VPWR VGND sg13g2_fill_2
X_3649_ _2053_ VPWR _2056_ VGND s0.was_valid_out\[2\][0] net967 sg13g2_o21ai_1
XFILLER_0_404 VPWR VGND sg13g2_fill_2
XFILLER_1_949 VPWR VGND sg13g2_decap_8
X_5319_ _0996_ _0997_ _0998_ VPWR VGND sg13g2_nor2_1
XFILLER_48_408 VPWR VGND sg13g2_decap_8
Xhold23 s0.was_valid_out\[3\][0] VPWR VGND net319 sg13g2_dlygate4sd3_1
XFILLER_0_459 VPWR VGND sg13g2_decap_8
Xhold12 s0.genblk1\[17\].modules.bubble VPWR VGND net308 sg13g2_dlygate4sd3_1
Xhold56 s0.data_out\[5\]\[5\] VPWR VGND net352 sg13g2_dlygate4sd3_1
Xhold45 s0.data_out\[17\]\[7\] VPWR VGND net341 sg13g2_dlygate4sd3_1
Xhold34 s0.data_out\[11\]\[4\] VPWR VGND net330 sg13g2_dlygate4sd3_1
XFILLER_29_56 VPWR VGND sg13g2_fill_2
Xhold67 s0.was_valid_out\[0\][0] VPWR VGND net363 sg13g2_dlygate4sd3_1
Xhold89 s0.data_out\[9\]\[5\] VPWR VGND net385 sg13g2_dlygate4sd3_1
Xhold78 s0.data_out\[0\]\[4\] VPWR VGND net374 sg13g2_dlygate4sd3_1
XFILLER_21_1004 VPWR VGND sg13g2_decap_8
XFILLER_17_839 VPWR VGND sg13g2_decap_8
XFILLER_16_316 VPWR VGND sg13g2_fill_2
XFILLER_29_699 VPWR VGND sg13g2_decap_8
XFILLER_12_511 VPWR VGND sg13g2_decap_8
XFILLER_24_371 VPWR VGND sg13g2_fill_2
XFILLER_25_894 VPWR VGND sg13g2_decap_8
XFILLER_12_522 VPWR VGND sg13g2_fill_1
XFILLER_8_515 VPWR VGND sg13g2_decap_8
XFILLER_8_559 VPWR VGND sg13g2_fill_1
Xfanout1010 net1011 net1010 VPWR VGND sg13g2_buf_2
Xfanout1021 net1022 net1021 VPWR VGND sg13g2_buf_8
XFILLER_48_920 VPWR VGND sg13g2_decap_8
Xfanout1032 net1034 net1032 VPWR VGND sg13g2_buf_8
Xfanout1043 net1044 net1043 VPWR VGND sg13g2_buf_8
X_6051__230 VPWR VGND net230 sg13g2_tiehi
XFILLER_0_971 VPWR VGND sg13g2_decap_8
Xfanout1054 net1056 net1054 VPWR VGND sg13g2_buf_2
Xfanout1065 net1068 net1065 VPWR VGND sg13g2_buf_8
Xfanout1098 net1099 net1098 VPWR VGND sg13g2_buf_8
Xfanout1076 net606 net1076 VPWR VGND sg13g2_buf_8
Xfanout1087 s0.valid_out\[10\][0] net1087 VPWR VGND sg13g2_buf_8
XFILLER_48_997 VPWR VGND sg13g2_decap_8
XFILLER_47_496 VPWR VGND sg13g2_decap_4
XFILLER_30_330 VPWR VGND sg13g2_fill_1
X_5670_ s0.data_out\[10\]\[7\] s0.data_out\[9\]\[7\] net1043 _1315_ VPWR VGND sg13g2_mux2_1
X_4621_ _0361_ net1155 _0320_ _0362_ VPWR VGND sg13g2_a21o_1
X_4552_ net1303 VPWR _0303_ VGND net406 _0298_ sg13g2_o21ai_1
X_3503_ VGND VPWR _1863_ _1921_ _1924_ net1253 sg13g2_a21oi_1
X_4483_ VGND VPWR net1168 s0.data_out\[18\]\[7\] _2800_ _2799_ sg13g2_a21oi_1
X_3434_ net993 VPWR _1859_ VGND _1857_ _1858_ sg13g2_o21ai_1
XFILLER_44_1004 VPWR VGND sg13g2_decap_8
X_3365_ _1797_ _1795_ _1798_ VPWR VGND _1796_ sg13g2_nand3b_1
X_6153_ net120 VGND VPWR _0203_ s0.data_out\[5\]\[1\] clknet_leaf_5_clk sg13g2_dfrbpq_2
X_5104_ net1115 net1060 _0801_ VPWR VGND sg13g2_nor2b_1
X_3296_ _1734_ net916 _1733_ VPWR VGND sg13g2_nand2_1
X_6084_ net194 VGND VPWR _0134_ s0.valid_out\[10\][0] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_5035_ _0738_ _0739_ _0737_ _0740_ VPWR VGND sg13g2_nand3_1
XFILLER_39_986 VPWR VGND sg13g2_decap_8
XFILLER_26_647 VPWR VGND sg13g2_decap_8
XFILLER_25_146 VPWR VGND sg13g2_decap_4
XFILLER_13_319 VPWR VGND sg13g2_fill_2
X_5937_ _1550_ VPWR _1551_ VGND _1543_ _1544_ sg13g2_o21ai_1
XFILLER_21_352 VPWR VGND sg13g2_decap_8
X_5868_ VGND VPWR _1489_ net526 net1328 sg13g2_or2_1
X_4819_ _0543_ net922 _0542_ VPWR VGND sg13g2_nand2_1
X_5799_ _1359_ VPWR _1425_ VGND net919 _1424_ sg13g2_o21ai_1
XFILLER_5_529 VPWR VGND sg13g2_decap_8
XFILLER_31_57 VPWR VGND sg13g2_decap_8
XFILLER_0_234 VPWR VGND sg13g2_fill_1
XFILLER_1_746 VPWR VGND sg13g2_decap_8
XFILLER_48_205 VPWR VGND sg13g2_decap_4
XFILLER_0_267 VPWR VGND sg13g2_fill_1
XFILLER_45_956 VPWR VGND sg13g2_decap_8
XFILLER_13_831 VPWR VGND sg13g2_fill_1
XFILLER_12_352 VPWR VGND sg13g2_decap_8
XFILLER_9_846 VPWR VGND sg13g2_fill_1
Xclkbuf_3_1__f_clk clknet_0_clk clknet_3_1__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_4_562 VPWR VGND sg13g2_fill_1
X_3150_ _1602_ net917 _1601_ VPWR VGND sg13g2_nand2_1
XFILLER_48_794 VPWR VGND sg13g2_decap_8
XFILLER_36_945 VPWR VGND sg13g2_decap_8
XFILLER_35_477 VPWR VGND sg13g2_fill_2
X_5722_ _1356_ _1357_ _0152_ VPWR VGND sg13g2_nor2_1
X_3983_ VGND VPWR net942 _2355_ _2356_ _2294_ sg13g2_a21oi_1
X_5653_ VGND VPWR _1298_ _1297_ net1270 sg13g2_or2_1
X_4604_ VGND VPWR _2829_ _0346_ _0347_ net1171 sg13g2_a21oi_1
XFILLER_30_193 VPWR VGND sg13g2_decap_4
X_5584_ _1237_ _1238_ _0133_ VPWR VGND sg13g2_nor2_1
Xhold301 s0.data_out\[13\]\[6\] VPWR VGND net597 sg13g2_dlygate4sd3_1
X_4535_ _2824_ _0273_ _0287_ _0288_ VPWR VGND sg13g2_or3_1
Xhold312 s0.data_out\[8\]\[2\] VPWR VGND net608 sg13g2_dlygate4sd3_1
X_4466_ net1170 net1053 _2785_ VPWR VGND sg13g2_nor2b_1
X_6205_ net27 VGND VPWR _0255_ s0.data_out\[1\]\[5\] clknet_leaf_9_clk sg13g2_dfrbpq_2
X_4397_ s0.data_out\[20\]\[5\] s0.data_out\[19\]\[5\] net1188 _2725_ VPWR VGND sg13g2_mux2_1
X_3417_ VGND VPWR net981 net533 _1844_ _1843_ sg13g2_a21oi_1
X_6136_ net139 VGND VPWR _0186_ s0.shift_out\[7\][0] clknet_leaf_17_clk sg13g2_dfrbpq_2
X_3348_ s0.data_out\[6\]\[3\] s0.data_out\[5\]\[3\] net999 _1781_ VPWR VGND sg13g2_mux2_1
X_6067_ net213 VGND VPWR _0117_ s0.data_out\[12\]\[6\] clknet_leaf_26_clk sg13g2_dfrbpq_2
X_3279_ _1719_ net463 net1008 VPWR VGND sg13g2_nand2b_1
X_5018_ s0.data_out\[15\]\[3\] s0.data_out\[14\]\[3\] net1130 _0723_ VPWR VGND sg13g2_mux2_1
XFILLER_27_956 VPWR VGND sg13g2_fill_1
XFILLER_42_915 VPWR VGND sg13g2_decap_8
XFILLER_26_79 VPWR VGND sg13g2_decap_8
XFILLER_13_127 VPWR VGND sg13g2_fill_1
XFILLER_13_149 VPWR VGND sg13g2_fill_1
XFILLER_22_650 VPWR VGND sg13g2_decap_8
XFILLER_42_78 VPWR VGND sg13g2_decap_8
XFILLER_10_878 VPWR VGND sg13g2_fill_2
XFILLER_1_543 VPWR VGND sg13g2_decap_8
XFILLER_49_569 VPWR VGND sg13g2_decap_8
XFILLER_18_901 VPWR VGND sg13g2_fill_1
XFILLER_45_753 VPWR VGND sg13g2_decap_8
XFILLER_44_263 VPWR VGND sg13g2_fill_2
XFILLER_13_650 VPWR VGND sg13g2_decap_4
XFILLER_5_860 VPWR VGND sg13g2_decap_8
X_4320_ VPWR _0017_ _2653_ VGND sg13g2_inv_1
X_4251_ _2591_ net1198 net523 VPWR VGND sg13g2_nand2_1
X_5996__290 VPWR VGND net290 sg13g2_tiehi
X_3202_ VGND VPWR _1648_ net517 net1329 sg13g2_or2_1
X_4182_ net1191 s0.data_out\[20\]\[2\] _2528_ VPWR VGND sg13g2_and2_1
X_3133_ net1005 _1584_ _1588_ VPWR VGND sg13g2_nor2_1
XFILLER_48_591 VPWR VGND sg13g2_decap_8
X_3966_ _2340_ net334 net956 VPWR VGND sg13g2_nand2b_1
X_5705_ net1061 net1260 net1224 _0147_ VPWR VGND sg13g2_mux2_1
X_3897_ VGND VPWR _2282_ net1208 net300 sg13g2_or2_1
X_5636_ net1039 net1051 _1283_ VPWR VGND sg13g2_nor2b_1
X_5567_ _1198_ _1210_ _1223_ _1224_ VPWR VGND sg13g2_or3_1
X_4518_ net1239 _2832_ _2834_ VPWR VGND sg13g2_nor2_1
Xhold142 s0.data_out\[15\]\[5\] VPWR VGND net438 sg13g2_dlygate4sd3_1
Xhold120 s0.data_out\[16\]\[4\] VPWR VGND net416 sg13g2_dlygate4sd3_1
X_5498_ _1158_ VPWR _1159_ VGND _1154_ _1157_ sg13g2_o21ai_1
Xhold153 _2297_ VPWR VGND net449 sg13g2_dlygate4sd3_1
Xhold131 _2189_ VPWR VGND net427 sg13g2_dlygate4sd3_1
Xhold186 s0.data_out\[8\]\[5\] VPWR VGND net482 sg13g2_dlygate4sd3_1
X_4449_ VGND VPWR _2703_ _2769_ _2770_ net1181 sg13g2_a21oi_1
Xhold175 s0.data_out\[13\]\[1\] VPWR VGND net471 sg13g2_dlygate4sd3_1
Xhold164 s0.data_out\[18\]\[0\] VPWR VGND net460 sg13g2_dlygate4sd3_1
Xhold197 s0.data_out\[18\]\[1\] VPWR VGND net493 sg13g2_dlygate4sd3_1
X_6119_ net157 VGND VPWR _0169_ s0.data_out\[8\]\[3\] clknet_leaf_15_clk sg13g2_dfrbpq_2
XFILLER_2_1001 VPWR VGND sg13g2_decap_8
XFILLER_27_742 VPWR VGND sg13g2_fill_2
XFILLER_27_753 VPWR VGND sg13g2_decap_8
XFILLER_42_778 VPWR VGND sg13g2_fill_2
XFILLER_23_992 VPWR VGND sg13g2_decap_8
XFILLER_5_112 VPWR VGND sg13g2_fill_2
XFILLER_5_134 VPWR VGND sg13g2_fill_1
XFILLER_49_311 VPWR VGND sg13g2_fill_2
XFILLER_2_896 VPWR VGND sg13g2_decap_8
XFILLER_49_366 VPWR VGND sg13g2_decap_8
XFILLER_49_344 VPWR VGND sg13g2_decap_4
XFILLER_18_753 VPWR VGND sg13g2_fill_1
XFILLER_45_550 VPWR VGND sg13g2_decap_8
XFILLER_45_583 VPWR VGND sg13g2_fill_2
XFILLER_32_222 VPWR VGND sg13g2_fill_2
XFILLER_33_723 VPWR VGND sg13g2_fill_1
X_3820_ _2205_ _2208_ net1298 _2209_ VPWR VGND sg13g2_nand3_1
XFILLER_32_266 VPWR VGND sg13g2_decap_4
X_3751_ s0.data_out\[3\]\[4\] s0.data_out\[2\]\[4\] net965 _2148_ VPWR VGND sg13g2_mux2_1
XFILLER_9_473 VPWR VGND sg13g2_fill_2
X_3682_ net960 net1064 _2084_ VPWR VGND sg13g2_nor2b_1
X_5421_ VGND VPWR net1105 _1089_ _1090_ _1049_ sg13g2_a21oi_1
X_5352_ VPWR _0113_ net505 VGND sg13g2_inv_1
X_4303_ _2638_ VPWR _2639_ VGND net1285 net462 sg13g2_o21ai_1
X_5283_ _0962_ _0963_ _0964_ VPWR VGND _0958_ sg13g2_nand3b_1
X_4234_ s0.data_out\[21\]\[1\] s0.data_out\[20\]\[1\] net1198 _2574_ VPWR VGND sg13g2_mux2_1
X_4165_ net1217 _2507_ _0002_ VPWR VGND sg13g2_nor2_1
X_3116_ _1573_ net1252 _1572_ VPWR VGND sg13g2_nand2_1
X_4096_ VPWR _2455_ net973 VGND sg13g2_inv_1
XFILLER_24_734 VPWR VGND sg13g2_fill_2
X_4998_ net1320 VPWR _0704_ VGND net921 _0703_ sg13g2_o21ai_1
X_3949_ VPWR _0254_ _2325_ VGND sg13g2_inv_1
X_5619_ _1268_ net934 _1267_ VPWR VGND sg13g2_nand2_1
XFILLER_47_815 VPWR VGND sg13g2_decap_8
XFILLER_48_44 VPWR VGND sg13g2_fill_2
XFILLER_27_561 VPWR VGND sg13g2_fill_2
XFILLER_42_531 VPWR VGND sg13g2_fill_1
XFILLER_14_233 VPWR VGND sg13g2_fill_1
XFILLER_42_597 VPWR VGND sg13g2_fill_1
XFILLER_9_38 VPWR VGND sg13g2_fill_1
XFILLER_30_737 VPWR VGND sg13g2_fill_2
XFILLER_31_1006 VPWR VGND sg13g2_decap_8
XFILLER_7_922 VPWR VGND sg13g2_decap_8
XFILLER_11_995 VPWR VGND sg13g2_decap_8
XFILLER_7_999 VPWR VGND sg13g2_decap_8
XFILLER_2_693 VPWR VGND sg13g2_decap_8
XFILLER_2_682 VPWR VGND sg13g2_decap_8
XFILLER_49_141 VPWR VGND sg13g2_fill_2
X_5993__293 VPWR VGND net293 sg13g2_tiehi
XFILLER_49_174 VPWR VGND sg13g2_decap_4
XFILLER_49_196 VPWR VGND sg13g2_decap_8
X_5970_ net46 VGND VPWR _0020_ s0.data_out\[20\]\[5\] clknet_leaf_2_clk sg13g2_dfrbpq_2
X_4921_ _0618_ _0620_ _0638_ VPWR VGND sg13g2_nor2b_1
X_4852_ net1137 s0.data_out\[15\]\[5\] _0572_ VPWR VGND sg13g2_and2_1
XFILLER_21_726 VPWR VGND sg13g2_fill_2
X_3803_ net1297 VPWR _2194_ VGND net930 _2193_ sg13g2_o21ai_1
X_6206__286 VPWR VGND net286 sg13g2_tiehi
X_4783_ s0.data_out\[17\]\[5\] s0.data_out\[16\]\[5\] net1154 _0512_ VPWR VGND sg13g2_mux2_1
X_3734_ s0.data_out\[3\]\[3\] s0.data_out\[2\]\[3\] net965 _2131_ VPWR VGND sg13g2_mux2_1
X_3665_ _2069_ net932 _2068_ VPWR VGND sg13g2_nand2_1
X_5404_ _1073_ net1102 _1072_ VPWR VGND sg13g2_nand2b_1
X_3596_ VGND VPWR net969 _2004_ _2005_ _1954_ sg13g2_a21oi_1
X_5335_ _1011_ VPWR _1012_ VGND net1335 net473 sg13g2_o21ai_1
X_5266_ _0903_ VPWR _0947_ VGND net935 _0946_ sg13g2_o21ai_1
X_4217_ net356 net1207 _2559_ VPWR VGND sg13g2_nor2b_1
X_5197_ VGND VPWR _2445_ _0882_ _0097_ _0887_ sg13g2_a21oi_1
X_4148_ s0.data_out\[21\]\[6\] net912 _2501_ VPWR VGND sg13g2_nor2_1
XFILLER_44_829 VPWR VGND sg13g2_decap_8
X_4079_ _2439_ VPWR _2440_ VGND _2436_ _2438_ sg13g2_o21ai_1
XFILLER_37_892 VPWR VGND sg13g2_fill_1
XFILLER_37_881 VPWR VGND sg13g2_fill_1
XFILLER_34_24 VPWR VGND sg13g2_decap_4
Xclkload1 clknet_3_7__leaf_clk clkload1/X VPWR VGND sg13g2_buf_8
XFILLER_4_914 VPWR VGND sg13g2_decap_8
Xfanout1203 net332 net1203 VPWR VGND sg13g2_buf_8
Xfanout1214 net1215 net1214 VPWR VGND sg13g2_buf_8
Xfanout1225 net1227 net1225 VPWR VGND sg13g2_buf_8
Xfanout1247 net1249 net1247 VPWR VGND sg13g2_buf_1
Xfanout1236 net1238 net1236 VPWR VGND sg13g2_buf_8
XFILLER_47_612 VPWR VGND sg13g2_decap_8
Xfanout1258 net1259 net1258 VPWR VGND sg13g2_buf_8
Xfanout1269 net1272 net1269 VPWR VGND sg13g2_buf_1
XFILLER_47_689 VPWR VGND sg13g2_decap_8
XFILLER_46_144 VPWR VGND sg13g2_decap_4
XFILLER_34_328 VPWR VGND sg13g2_fill_1
XFILLER_27_391 VPWR VGND sg13g2_fill_1
XFILLER_43_884 VPWR VGND sg13g2_decap_8
XFILLER_30_512 VPWR VGND sg13g2_decap_4
XFILLER_11_770 VPWR VGND sg13g2_fill_1
XFILLER_30_589 VPWR VGND sg13g2_fill_2
X_3450_ net1314 VPWR _1873_ VGND _2470_ _1872_ sg13g2_o21ai_1
X_3381_ _1795_ _1797_ _1814_ VPWR VGND sg13g2_nor2b_1
X_5120_ net1115 net1052 _0815_ VPWR VGND sg13g2_nor2b_1
X_5051_ _0741_ _0751_ _0728_ _0756_ VPWR VGND _0755_ sg13g2_nand4_1
X_4002_ _2375_ _2374_ net1241 _2371_ net1232 VPWR VGND sg13g2_a22oi_1
XFILLER_37_122 VPWR VGND sg13g2_fill_2
XFILLER_37_166 VPWR VGND sg13g2_fill_1
XFILLER_37_144 VPWR VGND sg13g2_fill_2
Xheichips25_top_sorter_21 VPWR VGND uio_out[6] sg13g2_tielo
Xheichips25_top_sorter_10 VPWR VGND uio_oe[0] sg13g2_tielo
XFILLER_37_177 VPWR VGND sg13g2_decap_8
XFILLER_25_339 VPWR VGND sg13g2_fill_2
X_5953_ net64 VGND VPWR net369 s0.data_out\[21\]\[0\] clknet_leaf_37_clk sg13g2_dfrbpq_1
X_4904_ _0620_ _0618_ _0621_ VPWR VGND _0619_ sg13g2_nand3b_1
X_5884_ _1499_ _1502_ net1328 _1503_ VPWR VGND sg13g2_nand3_1
X_4835_ VGND VPWR _0489_ _0556_ _0557_ net1149 sg13g2_a21oi_1
X_4766_ _0494_ VPWR _0495_ VGND _0487_ _0488_ sg13g2_o21ai_1
X_3717_ VGND VPWR _2115_ net515 net1309 sg13g2_or2_1
X_6177__94 VPWR VGND net94 sg13g2_tiehi
X_4697_ VGND VPWR _0433_ net496 net1304 sg13g2_or2_1
X_3648_ VPWR _2055_ _2054_ VGND sg13g2_inv_1
X_3579_ net1310 VPWR _1990_ VGND net914 _1989_ sg13g2_o21ai_1
XFILLER_1_928 VPWR VGND sg13g2_decap_8
X_5318_ net1229 net1098 _0997_ VPWR VGND sg13g2_nor2b_1
Xhold13 s0.genblk1\[6\].modules.bubble VPWR VGND net309 sg13g2_dlygate4sd3_1
XFILLER_0_438 VPWR VGND sg13g2_decap_8
Xhold24 _0224_ VPWR VGND net320 sg13g2_dlygate4sd3_1
Xhold46 _0471_ VPWR VGND net342 sg13g2_dlygate4sd3_1
X_5249_ net1107 net1052 _0932_ VPWR VGND sg13g2_nor2b_1
Xhold35 _1035_ VPWR VGND net331 sg13g2_dlygate4sd3_1
Xhold57 s0.was_valid_out\[4\][0] VPWR VGND net353 sg13g2_dlygate4sd3_1
Xhold68 s0.data_out\[21\]\[7\] VPWR VGND net364 sg13g2_dlygate4sd3_1
Xhold79 s0.was_valid_out\[17\][0] VPWR VGND net375 sg13g2_dlygate4sd3_1
XFILLER_29_656 VPWR VGND sg13g2_fill_1
XFILLER_45_12 VPWR VGND sg13g2_fill_1
XFILLER_43_147 VPWR VGND sg13g2_fill_1
Xfanout1011 s0.valid_out\[6\][0] net1011 VPWR VGND sg13g2_buf_8
Xfanout1022 s0.valid_out\[7\][0] net1022 VPWR VGND sg13g2_buf_8
XFILLER_0_950 VPWR VGND sg13g2_decap_8
Xfanout1000 net1003 net1000 VPWR VGND sg13g2_buf_8
Xfanout1055 net1056 net1055 VPWR VGND sg13g2_buf_8
Xfanout1033 net1034 net1033 VPWR VGND sg13g2_buf_2
Xfanout1044 s0.valid_out\[9\][0] net1044 VPWR VGND sg13g2_buf_2
Xfanout1088 net1090 net1088 VPWR VGND sg13g2_buf_8
Xfanout1066 net1068 net1066 VPWR VGND sg13g2_buf_8
Xfanout1077 net1078 net1077 VPWR VGND sg13g2_buf_8
XFILLER_48_976 VPWR VGND sg13g2_decap_8
XFILLER_47_442 VPWR VGND sg13g2_decap_8
Xfanout1099 net500 net1099 VPWR VGND sg13g2_buf_8
XFILLER_19_166 VPWR VGND sg13g2_decap_4
XFILLER_34_114 VPWR VGND sg13g2_decap_8
XFILLER_34_125 VPWR VGND sg13g2_fill_1
XFILLER_31_810 VPWR VGND sg13g2_fill_2
XFILLER_42_191 VPWR VGND sg13g2_decap_8
XFILLER_15_394 VPWR VGND sg13g2_decap_8
XFILLER_31_832 VPWR VGND sg13g2_fill_2
XFILLER_31_843 VPWR VGND sg13g2_fill_2
X_4620_ s0.data_out\[18\]\[2\] s0.data_out\[17\]\[2\] net1163 _0361_ VPWR VGND sg13g2_mux2_1
XFILLER_7_560 VPWR VGND sg13g2_decap_4
X_4551_ VGND VPWR _0296_ _0299_ _0302_ _0301_ sg13g2_a21oi_1
X_3502_ _1923_ _1922_ _1918_ VPWR VGND sg13g2_nand2b_1
X_4482_ net1168 net1045 _2799_ VPWR VGND sg13g2_nor2b_1
X_6221_ net71 VGND VPWR _0271_ s0.genblk1\[9\].modules.bubble clknet_leaf_18_clk sg13g2_dfrbpq_1
X_3433_ net982 net1058 _1858_ VPWR VGND sg13g2_nor2b_1
X_6152_ net121 VGND VPWR _0202_ s0.data_out\[5\]\[0\] clknet_leaf_5_clk sg13g2_dfrbpq_2
X_3364_ VGND VPWR _1797_ _1790_ net1235 sg13g2_or2_1
X_5103_ VGND VPWR _0742_ _0799_ _0800_ net1128 sg13g2_a21oi_1
XFILLER_32_0 VPWR VGND sg13g2_decap_8
X_3295_ s0.data_out\[5\]\[3\] s0.data_out\[6\]\[3\] net1008 _1733_ VPWR VGND sg13g2_mux2_1
X_6083_ net196 VGND VPWR net380 s0.was_valid_out\[10\][0] clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_38_420 VPWR VGND sg13g2_fill_1
X_5034_ VGND VPWR _0739_ _0736_ net1244 sg13g2_or2_1
XFILLER_39_965 VPWR VGND sg13g2_decap_8
XFILLER_13_309 VPWR VGND sg13g2_fill_1
XFILLER_15_48 VPWR VGND sg13g2_fill_2
X_5936_ _1550_ _1549_ net1266 _1535_ net1271 VPWR VGND sg13g2_a22oi_1
XFILLER_40_128 VPWR VGND sg13g2_decap_8
X_6028__255 VPWR VGND net255 sg13g2_tiehi
X_5867_ net1328 VPWR _1488_ VGND net918 _1487_ sg13g2_o21ai_1
X_4818_ s0.data_out\[15\]\[1\] s0.data_out\[16\]\[1\] net1152 _0542_ VPWR VGND sg13g2_mux2_1
XFILLER_21_397 VPWR VGND sg13g2_fill_1
X_5798_ VGND VPWR net1024 _1423_ _1424_ _1361_ sg13g2_a21oi_1
X_4749_ _0477_ net1144 _0437_ _0478_ VPWR VGND sg13g2_a21o_1
XFILLER_1_725 VPWR VGND sg13g2_decap_8
XFILLER_0_246 VPWR VGND sg13g2_decap_8
X_6215__149 VPWR VGND net149 sg13g2_tiehi
X_6035__248 VPWR VGND net248 sg13g2_tiehi
XFILLER_5_1021 VPWR VGND sg13g2_decap_8
XFILLER_29_420 VPWR VGND sg13g2_fill_1
XFILLER_29_442 VPWR VGND sg13g2_decap_8
XFILLER_45_935 VPWR VGND sg13g2_decap_8
XFILLER_16_114 VPWR VGND sg13g2_fill_2
XFILLER_17_615 VPWR VGND sg13g2_fill_2
XFILLER_17_637 VPWR VGND sg13g2_fill_1
XFILLER_16_136 VPWR VGND sg13g2_decap_8
XFILLER_24_191 VPWR VGND sg13g2_fill_2
XFILLER_8_324 VPWR VGND sg13g2_decap_4
XFILLER_12_364 VPWR VGND sg13g2_fill_1
XFILLER_4_596 VPWR VGND sg13g2_fill_1
XFILLER_48_773 VPWR VGND sg13g2_decap_8
XFILLER_35_456 VPWR VGND sg13g2_decap_8
XFILLER_22_106 VPWR VGND sg13g2_fill_2
X_3982_ s0.data_out\[1\]\[0\] s0.data_out\[0\]\[0\] net946 _2355_ VPWR VGND sg13g2_mux2_1
XFILLER_44_990 VPWR VGND sg13g2_decap_8
X_5721_ net1346 VPWR _1357_ VGND net453 _1352_ sg13g2_o21ai_1
X_5652_ VGND VPWR net1079 _1296_ _1297_ _1254_ sg13g2_a21oi_1
X_4603_ _0346_ s0.data_out\[17\]\[6\] net1177 VPWR VGND sg13g2_nand2b_1
X_5583_ net1344 VPWR _1238_ VGND net379 _1233_ sg13g2_o21ai_1
XFILLER_7_82 VPWR VGND sg13g2_decap_8
Xhold302 s0.data_out\[14\]\[6\] VPWR VGND net598 sg13g2_dlygate4sd3_1
X_4534_ _0282_ _0286_ _0278_ _0287_ VPWR VGND sg13g2_nand3_1
Xhold313 _1377_ VPWR VGND net609 sg13g2_dlygate4sd3_1
X_4465_ VGND VPWR _2724_ _2783_ _2784_ net1184 sg13g2_a21oi_1
X_4396_ _2724_ net1188 net586 VPWR VGND sg13g2_nand2_1
X_3416_ net981 net1066 _1843_ VPWR VGND sg13g2_nor2b_1
X_6204_ net40 VGND VPWR _0254_ s0.data_out\[1\]\[4\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_6135_ net140 VGND VPWR _0185_ s0.data_out\[7\]\[7\] clknet_leaf_17_clk sg13g2_dfrbpq_2
X_3347_ VPWR VGND _1713_ net1282 _1778_ net1277 _1780_ _1775_ sg13g2_a221oi_1
X_6066_ net214 VGND VPWR _0116_ s0.data_out\[12\]\[5\] clknet_leaf_26_clk sg13g2_dfrbpq_2
XFILLER_39_740 VPWR VGND sg13g2_fill_1
X_5017_ _0722_ net1271 _0666_ _0710_ VPWR VGND sg13g2_and3_1
X_3278_ VPWR _0190_ _1718_ VGND sg13g2_inv_1
XFILLER_26_36 VPWR VGND sg13g2_fill_1
XFILLER_26_434 VPWR VGND sg13g2_decap_8
XFILLER_41_415 VPWR VGND sg13g2_fill_1
XFILLER_42_24 VPWR VGND sg13g2_fill_2
XFILLER_42_13 VPWR VGND sg13g2_decap_8
X_5919_ s0.data_out\[8\]\[2\] s0.data_out\[7\]\[2\] net1019 _1533_ VPWR VGND sg13g2_mux2_1
XFILLER_10_824 VPWR VGND sg13g2_decap_8
XFILLER_6_828 VPWR VGND sg13g2_fill_2
XFILLER_10_857 VPWR VGND sg13g2_fill_2
X_6041__241 VPWR VGND net241 sg13g2_tiehi
XFILLER_1_522 VPWR VGND sg13g2_decap_8
XFILLER_49_548 VPWR VGND sg13g2_decap_8
XFILLER_1_599 VPWR VGND sg13g2_decap_8
XFILLER_45_732 VPWR VGND sg13g2_decap_8
XFILLER_44_220 VPWR VGND sg13g2_decap_8
XFILLER_17_423 VPWR VGND sg13g2_fill_1
XFILLER_33_916 VPWR VGND sg13g2_decap_4
XFILLER_32_426 VPWR VGND sg13g2_fill_2
XFILLER_41_982 VPWR VGND sg13g2_decap_8
XFILLER_12_172 VPWR VGND sg13g2_fill_1
XFILLER_34_1026 VPWR VGND sg13g2_fill_2
XFILLER_9_677 VPWR VGND sg13g2_fill_1
X_4250_ _2583_ _2589_ _2590_ VPWR VGND sg13g2_nor2_1
XFILLER_4_382 VPWR VGND sg13g2_decap_8
X_3201_ net1329 VPWR _1647_ VGND net917 _1646_ sg13g2_o21ai_1
X_4181_ VPWR _0004_ net371 VGND sg13g2_inv_1
X_3132_ _1586_ VPWR _1587_ VGND s0.was_valid_out\[6\][0] net1010 sg13g2_o21ai_1
XFILLER_48_570 VPWR VGND sg13g2_decap_8
X_3965_ VPWR _0256_ _2339_ VGND sg13g2_inv_1
X_3896_ _2170_ _2279_ _2280_ _2281_ VPWR VGND sg13g2_nor3_1
X_5704_ VGND VPWR net1223 net1211 _0146_ _1345_ sg13g2_a21oi_1
XFILLER_32_982 VPWR VGND sg13g2_decap_8
X_5635_ VGND VPWR _1203_ _1281_ _1282_ net1082 sg13g2_a21oi_1
X_6025__258 VPWR VGND net258 sg13g2_tiehi
XFILLER_12_49 VPWR VGND sg13g2_decap_8
Xhold110 s0.was_valid_out\[18\][0] VPWR VGND net406 sg13g2_dlygate4sd3_1
X_5566_ _1223_ _1218_ _1222_ VPWR VGND sg13g2_nand2_1
Xhold121 s0.data_out\[2\]\[4\] VPWR VGND net417 sg13g2_dlygate4sd3_1
Xhold143 s0.data_out\[13\]\[0\] VPWR VGND net439 sg13g2_dlygate4sd3_1
X_4517_ _2833_ _2832_ net1240 _2828_ net1231 VPWR VGND sg13g2_a22oi_1
Xhold132 s0.data_out\[9\]\[0\] VPWR VGND net428 sg13g2_dlygate4sd3_1
X_5497_ VGND VPWR _1158_ net330 net1337 sg13g2_or2_1
Xhold154 s0.data_out\[16\]\[0\] VPWR VGND net450 sg13g2_dlygate4sd3_1
X_4448_ _2769_ net478 net1187 VPWR VGND sg13g2_nand2b_1
Xhold165 s0.data_out\[15\]\[0\] VPWR VGND net461 sg13g2_dlygate4sd3_1
Xhold176 s0.data_out\[12\]\[3\] VPWR VGND net472 sg13g2_dlygate4sd3_1
Xhold187 _1518_ VPWR VGND net483 sg13g2_dlygate4sd3_1
Xhold198 _0317_ VPWR VGND net494 sg13g2_dlygate4sd3_1
X_4379_ _2707_ _2706_ net1260 _2691_ net1268 VPWR VGND sg13g2_a22oi_1
X_6118_ net158 VGND VPWR _0168_ s0.data_out\[8\]\[2\] clknet_leaf_22_clk sg13g2_dfrbpq_2
XFILLER_39_581 VPWR VGND sg13g2_fill_1
X_6049_ net232 VGND VPWR _0099_ s0.data_out\[13\]\[0\] clknet_leaf_29_clk sg13g2_dfrbpq_2
XFILLER_27_710 VPWR VGND sg13g2_decap_8
X_6205__27 VPWR VGND net27 sg13g2_tiehi
XFILLER_42_702 VPWR VGND sg13g2_fill_1
XFILLER_41_223 VPWR VGND sg13g2_fill_2
XFILLER_14_415 VPWR VGND sg13g2_fill_1
XFILLER_15_938 VPWR VGND sg13g2_fill_1
XFILLER_41_278 VPWR VGND sg13g2_fill_1
XFILLER_23_971 VPWR VGND sg13g2_decap_8
XFILLER_10_632 VPWR VGND sg13g2_fill_1
XFILLER_6_636 VPWR VGND sg13g2_fill_1
XFILLER_6_625 VPWR VGND sg13g2_decap_8
XFILLER_10_687 VPWR VGND sg13g2_fill_1
XFILLER_6_647 VPWR VGND sg13g2_fill_2
XFILLER_5_179 VPWR VGND sg13g2_fill_2
XFILLER_2_875 VPWR VGND sg13g2_decap_8
XFILLER_37_507 VPWR VGND sg13g2_decap_8
XFILLER_37_518 VPWR VGND sg13g2_fill_2
XFILLER_17_253 VPWR VGND sg13g2_decap_8
XFILLER_18_798 VPWR VGND sg13g2_fill_1
X_3750_ _2146_ _2144_ _2147_ VPWR VGND _2145_ sg13g2_nand3b_1
XFILLER_14_982 VPWR VGND sg13g2_decap_8
XFILLER_9_441 VPWR VGND sg13g2_decap_4
XFILLER_9_452 VPWR VGND sg13g2_decap_8
X_3681_ VGND VPWR _2013_ _2082_ _2083_ net971 sg13g2_a21oi_1
XFILLER_9_496 VPWR VGND sg13g2_fill_1
X_5420_ _1088_ net1091 _1050_ _1089_ VPWR VGND sg13g2_a21o_1
X_5351_ _1025_ VPWR _1026_ VGND _1021_ _1024_ sg13g2_o21ai_1
X_4302_ _2634_ _2637_ net1286 _2638_ VPWR VGND sg13g2_nand3_1
X_5282_ VGND VPWR _0963_ _0947_ net1212 sg13g2_or2_1
X_4233_ _2532_ VPWR _2573_ VGND _2457_ _2572_ sg13g2_o21ai_1
XFILLER_4_190 VPWR VGND sg13g2_fill_1
X_4164_ _2512_ _2513_ _0001_ VPWR VGND sg13g2_nor2_1
X_3115_ VGND VPWR net1026 _1571_ _1572_ _1513_ sg13g2_a21oi_1
X_4095_ VPWR _2454_ net1082 VGND sg13g2_inv_1
XFILLER_24_713 VPWR VGND sg13g2_fill_1
X_4997_ VGND VPWR net1123 s0.data_out\[14\]\[7\] _0703_ _0702_ sg13g2_a21oi_1
XFILLER_23_278 VPWR VGND sg13g2_fill_1
X_3948_ _2324_ VPWR _2325_ VGND net1298 net394 sg13g2_o21ai_1
X_3879_ VPWR _2264_ _2263_ VGND sg13g2_inv_1
X_5618_ s0.data_out\[9\]\[4\] s0.data_out\[10\]\[4\] net1086 _1267_ VPWR VGND sg13g2_mux2_1
XFILLER_3_617 VPWR VGND sg13g2_fill_2
X_5549_ VGND VPWR net1094 _1205_ _1206_ _1168_ sg13g2_a21oi_1
XFILLER_24_1014 VPWR VGND sg13g2_decap_8
XFILLER_9_17 VPWR VGND sg13g2_fill_1
XFILLER_23_790 VPWR VGND sg13g2_fill_2
XFILLER_11_974 VPWR VGND sg13g2_decap_8
XFILLER_10_484 VPWR VGND sg13g2_fill_1
XFILLER_7_978 VPWR VGND sg13g2_decap_8
XFILLER_36_7 VPWR VGND sg13g2_decap_4
XFILLER_2_661 VPWR VGND sg13g2_decap_8
X_4920_ _0621_ _0636_ _0637_ VPWR VGND sg13g2_nor2b_1
X_4851_ _0571_ net923 _0570_ VPWR VGND sg13g2_nand2_1
X_3802_ VGND VPWR net949 net458 _2193_ _2192_ sg13g2_a21oi_1
X_4782_ _0450_ VPWR _0511_ VGND net924 _0510_ sg13g2_o21ai_1
X_6189__81 VPWR VGND net81 sg13g2_tiehi
X_3733_ VPWR VGND _2128_ _2129_ _2124_ net1212 _2130_ _2120_ sg13g2_a221oi_1
X_3664_ s0.data_out\[2\]\[1\] s0.data_out\[3\]\[1\] net976 _2068_ VPWR VGND sg13g2_mux2_1
X_5403_ VGND VPWR net1088 _1071_ _1072_ _1009_ sg13g2_a21oi_1
X_3595_ s0.data_out\[4\]\[1\] s0.data_out\[3\]\[1\] net976 _2004_ VPWR VGND sg13g2_mux2_1
XFILLER_47_1025 VPWR VGND sg13g2_decap_4
X_5334_ _1007_ _1010_ net1335 _1011_ VPWR VGND sg13g2_nand3_1
X_5265_ VGND VPWR net1101 _0945_ _0946_ _0905_ sg13g2_a21oi_1
X_5196_ net1338 VPWR _0887_ VGND _0884_ _0886_ sg13g2_o21ai_1
X_4216_ net1204 VPWR _2558_ VGND _2556_ _2557_ sg13g2_o21ai_1
XFILLER_18_26 VPWR VGND sg13g2_decap_8
X_4147_ _2500_ VPWR net7 VGND _2475_ net912 sg13g2_o21ai_1
XFILLER_29_816 VPWR VGND sg13g2_fill_1
XFILLER_44_808 VPWR VGND sg13g2_decap_8
X_4078_ VGND VPWR net1232 _2425_ _2439_ net1227 sg13g2_a21oi_1
XFILLER_34_58 VPWR VGND sg13g2_fill_2
XFILLER_24_598 VPWR VGND sg13g2_decap_8
XFILLER_7_219 VPWR VGND sg13g2_fill_2
XFILLER_7_208 VPWR VGND sg13g2_decap_8
Xclkload2 VPWR clkload2/Y clknet_leaf_0_clk VGND sg13g2_inv_1
XFILLER_11_259 VPWR VGND sg13g2_fill_2
XFILLER_1_4 VPWR VGND sg13g2_decap_8
Xfanout1204 net332 net1204 VPWR VGND sg13g2_buf_8
Xfanout1226 net1227 net1226 VPWR VGND sg13g2_buf_8
Xfanout1237 net1238 net1237 VPWR VGND sg13g2_buf_8
Xfanout1215 _2476_ net1215 VPWR VGND sg13g2_buf_8
XFILLER_47_602 VPWR VGND sg13g2_decap_4
Xfanout1259 ui_in[4] net1259 VPWR VGND sg13g2_buf_8
Xfanout1248 net1249 net1248 VPWR VGND sg13g2_buf_8
XFILLER_46_101 VPWR VGND sg13g2_decap_4
XFILLER_47_668 VPWR VGND sg13g2_decap_8
XFILLER_27_370 VPWR VGND sg13g2_fill_2
XFILLER_28_893 VPWR VGND sg13g2_fill_1
XFILLER_43_863 VPWR VGND sg13g2_decap_8
XFILLER_7_742 VPWR VGND sg13g2_fill_2
XFILLER_7_775 VPWR VGND sg13g2_decap_8
X_3380_ _1798_ _1812_ _1813_ VPWR VGND sg13g2_nor2b_1
XFILLER_3_992 VPWR VGND sg13g2_decap_8
X_5050_ _0752_ _0753_ _0754_ _0755_ VPWR VGND sg13g2_nor3_1
X_4001_ VGND VPWR net952 _2373_ _2374_ _2334_ sg13g2_a21oi_1
Xheichips25_top_sorter_22 VPWR VGND uio_out[7] sg13g2_tielo
Xheichips25_top_sorter_11 VPWR VGND uio_oe[1] sg13g2_tielo
X_5952_ net65 VGND VPWR _0002_ s0.valid_out\[21\][0] clknet_leaf_2_clk sg13g2_dfrbpq_2
X_4903_ VGND VPWR _0620_ _0613_ net1235 sg13g2_or2_1
X_5883_ net1023 VPWR _1502_ VGND _1500_ _1501_ sg13g2_o21ai_1
X_4834_ _0556_ net387 net1152 VPWR VGND sg13g2_nand2b_1
XFILLER_21_535 VPWR VGND sg13g2_fill_1
X_4765_ _0494_ _0493_ net1262 _0479_ net1268 VPWR VGND sg13g2_a22oi_1
XFILLER_14_1024 VPWR VGND sg13g2_decap_4
X_3716_ net1309 VPWR _2114_ VGND net933 _2113_ sg13g2_o21ai_1
X_4696_ net1304 VPWR _0432_ VGND net924 _0431_ sg13g2_o21ai_1
X_3647_ VGND VPWR net932 _1935_ _2054_ _2053_ sg13g2_a21oi_1
XFILLER_20_38 VPWR VGND sg13g2_decap_4
X_3578_ VGND VPWR net972 s0.data_out\[3\]\[6\] _1989_ _1988_ sg13g2_a21oi_1
XFILLER_1_907 VPWR VGND sg13g2_decap_8
XFILLER_0_417 VPWR VGND sg13g2_decap_8
X_5317_ net1106 VPWR _0996_ VGND net1092 net1229 sg13g2_o21ai_1
Xhold14 s0.genblk1\[16\].modules.bubble VPWR VGND net310 sg13g2_dlygate4sd3_1
Xhold47 s0.shift_out\[9\][0] VPWR VGND net343 sg13g2_dlygate4sd3_1
X_5248_ VGND VPWR _0850_ _0930_ _0931_ net1117 sg13g2_a21oi_1
Xhold25 s0.was_valid_out\[16\][0] VPWR VGND net321 sg13g2_dlygate4sd3_1
Xhold36 s0.shift_out\[21\][0] VPWR VGND net332 sg13g2_dlygate4sd3_1
XFILLER_29_58 VPWR VGND sg13g2_fill_1
Xhold58 s0.shift_out\[0\][0] VPWR VGND net354 sg13g2_dlygate4sd3_1
X_5179_ _0845_ _0857_ _0869_ _0871_ _0872_ VPWR VGND sg13g2_or4_1
Xhold69 _0010_ VPWR VGND net365 sg13g2_dlygate4sd3_1
XFILLER_17_808 VPWR VGND sg13g2_decap_8
XFILLER_44_649 VPWR VGND sg13g2_fill_1
XFILLER_44_638 VPWR VGND sg13g2_fill_2
XFILLER_45_57 VPWR VGND sg13g2_fill_2
XFILLER_24_373 VPWR VGND sg13g2_fill_1
XFILLER_12_568 VPWR VGND sg13g2_fill_2
XFILLER_4_723 VPWR VGND sg13g2_fill_2
Xfanout1001 net1002 net1001 VPWR VGND sg13g2_buf_2
Xfanout1012 net340 net1012 VPWR VGND sg13g2_buf_8
Xfanout1034 s0.valid_out\[8\][0] net1034 VPWR VGND sg13g2_buf_8
Xfanout1045 net1048 net1045 VPWR VGND sg13g2_buf_8
Xfanout1056 net607 net1056 VPWR VGND sg13g2_buf_8
Xfanout1023 net1026 net1023 VPWR VGND sg13g2_buf_8
XFILLER_48_955 VPWR VGND sg13g2_decap_8
XFILLER_47_421 VPWR VGND sg13g2_decap_4
Xfanout1089 net1090 net1089 VPWR VGND sg13g2_buf_1
Xfanout1067 net1068 net1067 VPWR VGND sg13g2_buf_1
Xfanout1078 net1079 net1078 VPWR VGND sg13g2_buf_8
XFILLER_43_660 VPWR VGND sg13g2_decap_8
XFILLER_37_1013 VPWR VGND sg13g2_decap_8
XFILLER_34_159 VPWR VGND sg13g2_decap_8
XFILLER_15_373 VPWR VGND sg13g2_fill_2
XFILLER_30_321 VPWR VGND sg13g2_fill_2
XFILLER_35_90 VPWR VGND sg13g2_fill_1
X_4550_ _0300_ VPWR _0301_ VGND net1158 _0294_ sg13g2_o21ai_1
X_3501_ _1863_ _1921_ net1253 _1922_ VPWR VGND sg13g2_nand3_1
XFILLER_7_594 VPWR VGND sg13g2_fill_1
X_4481_ VGND VPWR _2709_ _2797_ _2798_ net1185 sg13g2_a21oi_1
X_6220_ net84 VGND VPWR _0270_ s0.shift_out\[0\][0] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_6174__98 VPWR VGND net98 sg13g2_tiehi
X_3432_ net982 s0.data_out\[4\]\[4\] _1857_ VPWR VGND sg13g2_and2_1
X_6151_ net122 VGND VPWR _0201_ s0.valid_out\[5\][0] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_3363_ net1244 _1794_ _1796_ VPWR VGND sg13g2_nor2_1
X_5102_ _0799_ net430 net1132 VPWR VGND sg13g2_nand2b_1
X_6082_ net197 VGND VPWR _0132_ s0.genblk1\[10\].modules.bubble clknet_leaf_19_clk
+ sg13g2_dfrbpq_1
X_3294_ VPWR _0192_ net485 VGND sg13g2_inv_1
XFILLER_39_944 VPWR VGND sg13g2_decap_8
X_5033_ VGND VPWR _0738_ _0732_ net1235 sg13g2_or2_1
XFILLER_38_476 VPWR VGND sg13g2_fill_1
X_6167__105 VPWR VGND net105 sg13g2_tiehi
XFILLER_40_107 VPWR VGND sg13g2_decap_8
X_5935_ _1499_ _1548_ _1549_ VPWR VGND sg13g2_and2_1
XFILLER_34_671 VPWR VGND sg13g2_fill_2
XFILLER_22_822 VPWR VGND sg13g2_fill_2
X_5866_ VGND VPWR net1013 net419 _1487_ _1486_ sg13g2_a21oi_1
X_4817_ VPWR _0063_ _0541_ VGND sg13g2_inv_1
X_5797_ s0.data_out\[9\]\[0\] s0.data_out\[8\]\[0\] net1031 _1423_ VPWR VGND sg13g2_mux2_1
X_4748_ s0.data_out\[17\]\[2\] s0.data_out\[16\]\[2\] net1151 _0477_ VPWR VGND sg13g2_mux2_1
X_4679_ _0416_ _0417_ _0418_ VPWR VGND sg13g2_nor2b_1
XFILLER_1_704 VPWR VGND sg13g2_decap_8
XFILLER_5_1000 VPWR VGND sg13g2_decap_8
XFILLER_45_914 VPWR VGND sg13g2_decap_8
XFILLER_16_104 VPWR VGND sg13g2_decap_4
XFILLER_17_649 VPWR VGND sg13g2_fill_1
XFILLER_48_752 VPWR VGND sg13g2_decap_8
XFILLER_47_251 VPWR VGND sg13g2_decap_4
XFILLER_35_402 VPWR VGND sg13g2_fill_1
X_3981_ _2299_ _2353_ net1274 _2354_ VPWR VGND sg13g2_nand3_1
X_5720_ VGND VPWR _1350_ _1353_ _1356_ _1355_ sg13g2_a21oi_1
X_5651_ _1295_ net1040 _1255_ _1296_ VPWR VGND sg13g2_a21o_1
XFILLER_31_696 VPWR VGND sg13g2_fill_2
X_4602_ VPWR _0044_ net571 VGND sg13g2_inv_1
X_5582_ VGND VPWR _1231_ _1234_ _1237_ _1236_ sg13g2_a21oi_1
XFILLER_11_1016 VPWR VGND sg13g2_decap_8
XFILLER_11_1027 VPWR VGND sg13g2_fill_2
X_4533_ _0283_ _0284_ _0285_ _0286_ VPWR VGND sg13g2_nor3_1
Xhold314 s0.data_out\[8\]\[5\] VPWR VGND net610 sg13g2_dlygate4sd3_1
Xhold303 s0.data_out\[13\]\[5\] VPWR VGND net599 sg13g2_dlygate4sd3_1
X_4464_ _2783_ net570 net1189 VPWR VGND sg13g2_nand2b_1
X_6203_ net53 VGND VPWR _0253_ s0.data_out\[1\]\[3\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_4395_ _2662_ VPWR _2723_ VGND net931 _2722_ sg13g2_o21ai_1
X_3415_ VGND VPWR _1768_ _1841_ _1842_ net990 sg13g2_a21oi_1
X_6134_ net141 VGND VPWR _0184_ s0.data_out\[7\]\[6\] clknet_leaf_17_clk sg13g2_dfrbpq_2
X_3346_ _1772_ VPWR _1779_ VGND net1277 _1775_ sg13g2_o21ai_1
X_6065_ net215 VGND VPWR _0115_ s0.data_out\[12\]\[4\] clknet_leaf_26_clk sg13g2_dfrbpq_2
X_5016_ _0711_ VPWR _0721_ VGND net1277 _0716_ sg13g2_o21ai_1
X_3277_ _1717_ VPWR _1718_ VGND net1326 net412 sg13g2_o21ai_1
XFILLER_39_796 VPWR VGND sg13g2_fill_1
XFILLER_39_774 VPWR VGND sg13g2_fill_2
XFILLER_26_15 VPWR VGND sg13g2_decap_8
XFILLER_26_413 VPWR VGND sg13g2_fill_2
XFILLER_27_925 VPWR VGND sg13g2_fill_1
XFILLER_26_479 VPWR VGND sg13g2_fill_1
X_5918_ VPWR _0173_ net596 VGND sg13g2_inv_1
Xclkbuf_leaf_33_clk clknet_3_1__leaf_clk clknet_leaf_33_clk VPWR VGND sg13g2_buf_8
X_5849_ net1016 _1468_ _1473_ VPWR VGND sg13g2_nor2_1
XFILLER_1_578 VPWR VGND sg13g2_decap_8
XFILLER_27_1023 VPWR VGND sg13g2_decap_4
XFILLER_49_527 VPWR VGND sg13g2_decap_8
XFILLER_45_711 VPWR VGND sg13g2_decap_8
XFILLER_45_788 VPWR VGND sg13g2_decap_8
XFILLER_26_980 VPWR VGND sg13g2_decap_8
XFILLER_41_961 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_24_clk clknet_3_4__leaf_clk clknet_leaf_24_clk VPWR VGND sg13g2_buf_8
XFILLER_34_1005 VPWR VGND sg13g2_decap_8
XFILLER_13_674 VPWR VGND sg13g2_decap_8
XFILLER_8_144 VPWR VGND sg13g2_fill_2
XFILLER_5_895 VPWR VGND sg13g2_decap_8
X_3200_ VGND VPWR net1006 s0.data_out\[6\]\[7\] _1646_ _1645_ sg13g2_a21oi_1
X_4180_ _2526_ VPWR _2527_ VGND net1285 net370 sg13g2_o21ai_1
X_3131_ _1584_ _1585_ _1586_ VPWR VGND sg13g2_nor2_1
X_6018__266 VPWR VGND net266 sg13g2_tiehi
XFILLER_36_755 VPWR VGND sg13g2_decap_4
XFILLER_35_221 VPWR VGND sg13g2_fill_1
XFILLER_24_917 VPWR VGND sg13g2_fill_1
X_6164__108 VPWR VGND net108 sg13g2_tiehi
XFILLER_17_991 VPWR VGND sg13g2_decap_8
X_3964_ _2338_ VPWR _2339_ VGND _2334_ _2337_ sg13g2_o21ai_1
Xclkbuf_leaf_15_clk clknet_3_6__leaf_clk clknet_leaf_15_clk VPWR VGND sg13g2_buf_8
XFILLER_32_961 VPWR VGND sg13g2_decap_8
X_3895_ _2260_ _2261_ _2280_ VPWR VGND sg13g2_nor2b_1
X_5703_ net1224 net1065 _1345_ VPWR VGND sg13g2_nor2_1
X_5634_ _1281_ s0.data_out\[9\]\[6\] net1086 VPWR VGND sg13g2_nand2b_1
X_5565_ _1219_ _1220_ _1221_ _1222_ VPWR VGND sg13g2_nor3_1
Xhold100 s0.data_out\[1\]\[1\] VPWR VGND net396 sg13g2_dlygate4sd3_1
X_4516_ VGND VPWR net1184 _2831_ _2832_ _2791_ sg13g2_a21oi_1
Xhold111 _0037_ VPWR VGND net407 sg13g2_dlygate4sd3_1
Xhold144 s0.data_out\[4\]\[0\] VPWR VGND net440 sg13g2_dlygate4sd3_1
X_5496_ net1337 VPWR _1157_ VGND net939 _1156_ sg13g2_o21ai_1
Xhold122 s0.data_out\[10\]\[1\] VPWR VGND net418 sg13g2_dlygate4sd3_1
Xhold133 s0.data_out\[10\]\[4\] VPWR VGND net429 sg13g2_dlygate4sd3_1
X_4447_ VPWR _0029_ _2768_ VGND sg13g2_inv_1
Xhold166 s0.data_out\[20\]\[0\] VPWR VGND net462 sg13g2_dlygate4sd3_1
Xhold177 s0.data_out\[12\]\[0\] VPWR VGND net473 sg13g2_dlygate4sd3_1
Xhold155 s0.data_out\[9\]\[2\] VPWR VGND net451 sg13g2_dlygate4sd3_1
Xhold199 s0.data_out\[1\]\[7\] VPWR VGND net495 sg13g2_dlygate4sd3_1
Xhold188 s0.data_out\[6\]\[2\] VPWR VGND net484 sg13g2_dlygate4sd3_1
X_4378_ VGND VPWR net1193 _2705_ _2706_ _2655_ sg13g2_a21oi_1
X_6117_ net159 VGND VPWR _0167_ s0.data_out\[8\]\[1\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_3329_ net996 net1047 _1763_ VPWR VGND sg13g2_nor2b_1
XFILLER_37_36 VPWR VGND sg13g2_fill_2
X_6048_ net233 VGND VPWR _0098_ s0.valid_out\[13\][0] clknet_leaf_27_clk sg13g2_dfrbpq_2
XFILLER_37_69 VPWR VGND sg13g2_fill_2
XFILLER_27_744 VPWR VGND sg13g2_fill_1
XFILLER_26_254 VPWR VGND sg13g2_fill_1
XFILLER_26_287 VPWR VGND sg13g2_decap_4
XFILLER_23_950 VPWR VGND sg13g2_decap_8
XFILLER_30_909 VPWR VGND sg13g2_fill_2
XFILLER_10_655 VPWR VGND sg13g2_fill_2
XFILLER_6_659 VPWR VGND sg13g2_decap_8
XFILLER_5_114 VPWR VGND sg13g2_fill_1
XFILLER_5_147 VPWR VGND sg13g2_decap_8
XFILLER_2_854 VPWR VGND sg13g2_decap_8
XFILLER_49_313 VPWR VGND sg13g2_fill_1
XFILLER_45_585 VPWR VGND sg13g2_fill_1
XFILLER_21_909 VPWR VGND sg13g2_decap_4
XFILLER_14_961 VPWR VGND sg13g2_decap_8
XFILLER_43_90 VPWR VGND sg13g2_decap_4
XFILLER_9_420 VPWR VGND sg13g2_decap_8
XFILLER_40_290 VPWR VGND sg13g2_decap_8
X_3680_ _2082_ net446 net976 VPWR VGND sg13g2_nand2b_1
X_5350_ VGND VPWR _1025_ net504 net1332 sg13g2_or2_1
X_4301_ net1193 VPWR _2637_ VGND _2635_ _2636_ sg13g2_o21ai_1
X_5281_ _0962_ net1265 _0961_ VPWR VGND sg13g2_nand2_1
X_4232_ VGND VPWR net1191 _2571_ _2572_ _2529_ sg13g2_a21oi_1
Xclkbuf_leaf_4_clk clknet_3_1__leaf_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
X_4163_ net1291 VPWR _2513_ VGND net372 _2507_ sg13g2_o21ai_1
X_3114_ _1570_ net1016 _1514_ _1571_ VPWR VGND sg13g2_a21o_1
X_4094_ VPWR _2453_ net1118 VGND sg13g2_inv_1
XFILLER_49_891 VPWR VGND sg13g2_decap_8
X_6031__252 VPWR VGND net252 sg13g2_tiehi
XFILLER_24_736 VPWR VGND sg13g2_fill_1
X_4996_ net1123 net1047 _0702_ VPWR VGND sg13g2_nor2b_1
XFILLER_23_224 VPWR VGND sg13g2_fill_2
X_3947_ _2320_ _2323_ net1298 _2324_ VPWR VGND sg13g2_nand3_1
XFILLER_20_920 VPWR VGND sg13g2_decap_4
X_3878_ _2261_ _2262_ _2260_ _2263_ VPWR VGND sg13g2_nand3_1
XFILLER_20_997 VPWR VGND sg13g2_decap_8
X_5617_ VPWR _0138_ _1266_ VGND sg13g2_inv_1
X_6099__179 VPWR VGND net179 sg13g2_tiehi
X_5548_ _1204_ net1081 _1169_ _1205_ VPWR VGND sg13g2_a21o_1
X_5479_ VGND VPWR net1078 net506 _1142_ _1141_ sg13g2_a21oi_1
XFILLER_48_46 VPWR VGND sg13g2_fill_1
XFILLER_48_35 VPWR VGND sg13g2_decap_4
XFILLER_27_585 VPWR VGND sg13g2_decap_8
XFILLER_42_555 VPWR VGND sg13g2_fill_2
XFILLER_14_224 VPWR VGND sg13g2_fill_2
XFILLER_30_739 VPWR VGND sg13g2_fill_1
XFILLER_11_953 VPWR VGND sg13g2_decap_8
XFILLER_7_957 VPWR VGND sg13g2_decap_8
XFILLER_6_478 VPWR VGND sg13g2_fill_2
X_6015__269 VPWR VGND net269 sg13g2_tiehi
Xclkbuf_3_7__f_clk clknet_0_clk clknet_3_7__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_46_894 VPWR VGND sg13g2_decap_8
X_4850_ s0.data_out\[15\]\[5\] s0.data_out\[16\]\[5\] net1153 _0570_ VPWR VGND sg13g2_mux2_1
XFILLER_33_544 VPWR VGND sg13g2_decap_8
XFILLER_21_728 VPWR VGND sg13g2_fill_1
X_3801_ net949 net1065 _2192_ VPWR VGND sg13g2_nor2b_1
XFILLER_33_566 VPWR VGND sg13g2_decap_4
X_4781_ VGND VPWR net1146 _0509_ _0510_ _0452_ sg13g2_a21oi_1
XFILLER_20_249 VPWR VGND sg13g2_decap_8
X_3732_ VGND VPWR _2069_ _2123_ _2129_ net1276 sg13g2_a21oi_1
X_3663_ VPWR _0226_ _2067_ VGND sg13g2_inv_1
X_5402_ s0.data_out\[12\]\[0\] s0.data_out\[11\]\[0\] net1096 _1071_ VPWR VGND sg13g2_mux2_1
XFILLER_47_1004 VPWR VGND sg13g2_decap_8
X_5333_ net1102 VPWR _1010_ VGND _1008_ _1009_ sg13g2_o21ai_1
X_3594_ VGND VPWR _2003_ _2002_ net1269 sg13g2_or2_1
X_5264_ _0944_ VPWR _0945_ VGND net1108 _2487_ sg13g2_o21ai_1
X_5195_ _0886_ _0883_ _0885_ VPWR VGND sg13g2_nand2_1
X_4215_ net1195 net1049 _2557_ VPWR VGND sg13g2_nor2b_1
X_4146_ _2500_ net1246 net912 VPWR VGND sg13g2_nand2_1
XFILLER_18_38 VPWR VGND sg13g2_fill_2
X_4077_ _2437_ VPWR _2438_ VGND net1232 _2425_ sg13g2_o21ai_1
XFILLER_34_48 VPWR VGND sg13g2_fill_1
X_4979_ _0687_ _2464_ _0686_ VPWR VGND sg13g2_nand2_1
Xclkload3 VPWR clkload3/Y clknet_leaf_2_clk VGND sg13g2_inv_1
XFILLER_20_783 VPWR VGND sg13g2_decap_4
XFILLER_4_949 VPWR VGND sg13g2_decap_8
Xfanout1205 net332 net1205 VPWR VGND sg13g2_buf_1
Xfanout1227 uio_in[0] net1227 VPWR VGND sg13g2_buf_8
Xfanout1238 ui_in[7] net1238 VPWR VGND sg13g2_buf_8
XFILLER_8_1020 VPWR VGND sg13g2_decap_8
Xfanout1216 net1218 net1216 VPWR VGND sg13g2_buf_8
Xfanout1249 ui_in[5] net1249 VPWR VGND sg13g2_buf_8
XFILLER_47_647 VPWR VGND sg13g2_decap_8
XFILLER_35_809 VPWR VGND sg13g2_decap_8
XFILLER_28_861 VPWR VGND sg13g2_fill_1
XFILLER_43_842 VPWR VGND sg13g2_decap_8
XFILLER_27_382 VPWR VGND sg13g2_decap_8
XFILLER_11_761 VPWR VGND sg13g2_decap_8
X_6186__85 VPWR VGND net85 sg13g2_tiehi
XFILLER_10_260 VPWR VGND sg13g2_decap_4
XFILLER_6_253 VPWR VGND sg13g2_decap_8
XFILLER_6_286 VPWR VGND sg13g2_fill_1
XFILLER_3_971 VPWR VGND sg13g2_decap_8
XFILLER_2_481 VPWR VGND sg13g2_fill_2
X_4000_ _2372_ net943 _2335_ _2373_ VPWR VGND sg13g2_a21o_1
XFILLER_27_4 VPWR VGND sg13g2_fill_2
XFILLER_37_102 VPWR VGND sg13g2_fill_2
Xheichips25_top_sorter_12 VPWR VGND uio_oe[3] sg13g2_tielo
X_5951_ net67 VGND VPWR net373 s0.was_valid_out\[21\][0] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_6089__189 VPWR VGND net189 sg13g2_tiehi
XFILLER_34_820 VPWR VGND sg13g2_fill_2
XFILLER_46_691 VPWR VGND sg13g2_decap_8
X_4902_ net1244 _0617_ _0619_ VPWR VGND sg13g2_nor2_1
XFILLER_33_330 VPWR VGND sg13g2_fill_1
X_5882_ net1014 net1063 _1501_ VPWR VGND sg13g2_nor2b_1
X_4833_ VPWR _0065_ _0555_ VGND sg13g2_inv_1
X_4764_ _0443_ _0492_ _0493_ VPWR VGND sg13g2_and2_1
XFILLER_14_1003 VPWR VGND sg13g2_decap_8
X_3715_ VGND VPWR net963 s0.data_out\[2\]\[7\] _2113_ _2112_ sg13g2_a21oi_1
X_4695_ VGND VPWR net1144 net476 _0431_ _0430_ sg13g2_a21oi_1
X_3646_ _2051_ _2052_ _2053_ VPWR VGND sg13g2_nor2_1
X_3577_ net974 net1050 _1988_ VPWR VGND sg13g2_nor2b_1
X_5316_ net1337 net302 _0108_ VPWR VGND sg13g2_and2_1
X_5247_ _0930_ net588 net1121 VPWR VGND sg13g2_nand2b_1
Xhold15 s0.genblk1\[3\].modules.bubble VPWR VGND net311 sg13g2_dlygate4sd3_1
Xhold37 s0.shift_out\[20\][0] VPWR VGND net333 sg13g2_dlygate4sd3_1
Xhold26 _0061_ VPWR VGND net322 sg13g2_dlygate4sd3_1
Xhold59 s0.data_out\[3\]\[5\] VPWR VGND net355 sg13g2_dlygate4sd3_1
Xhold48 s0.data_out\[0\]\[5\] VPWR VGND net344 sg13g2_dlygate4sd3_1
X_5178_ _0867_ _0870_ _0861_ _0871_ VPWR VGND sg13g2_nand3_1
XFILLER_21_1018 VPWR VGND sg13g2_decap_8
X_4129_ VPWR _2488_ s0.data_out\[12\]\[3\] VGND sg13g2_inv_1
XFILLER_40_812 VPWR VGND sg13g2_fill_1
XFILLER_36_190 VPWR VGND sg13g2_fill_2
XFILLER_25_864 VPWR VGND sg13g2_fill_2
XFILLER_40_856 VPWR VGND sg13g2_fill_1
XFILLER_8_529 VPWR VGND sg13g2_fill_2
XFILLER_20_580 VPWR VGND sg13g2_fill_2
XFILLER_20_591 VPWR VGND sg13g2_fill_1
X_6183__88 VPWR VGND net88 sg13g2_tiehi
XFILLER_4_768 VPWR VGND sg13g2_decap_8
XFILLER_3_234 VPWR VGND sg13g2_fill_1
XFILLER_4_779 VPWR VGND sg13g2_fill_2
Xfanout1013 net1014 net1013 VPWR VGND sg13g2_buf_2
Xfanout1002 net1003 net1002 VPWR VGND sg13g2_buf_1
Xfanout1046 net1048 net1046 VPWR VGND sg13g2_buf_8
Xfanout1024 net1026 net1024 VPWR VGND sg13g2_buf_1
Xfanout1035 net1036 net1035 VPWR VGND sg13g2_buf_8
XFILLER_48_934 VPWR VGND sg13g2_decap_8
XFILLER_0_985 VPWR VGND sg13g2_decap_8
Xfanout1068 net600 net1068 VPWR VGND sg13g2_buf_8
Xfanout1057 net1060 net1057 VPWR VGND sg13g2_buf_8
Xfanout1079 net358 net1079 VPWR VGND sg13g2_buf_8
XFILLER_19_92 VPWR VGND sg13g2_decap_8
XFILLER_35_617 VPWR VGND sg13g2_fill_2
XFILLER_15_352 VPWR VGND sg13g2_fill_2
X_3500_ _1921_ net994 _1920_ VPWR VGND sg13g2_nand2b_1
X_4480_ _2797_ s0.data_out\[18\]\[7\] net1187 VPWR VGND sg13g2_nand2b_1
X_3431_ _1856_ net915 _1855_ VPWR VGND sg13g2_nand2_1
X_6150_ net124 VGND VPWR net384 s0.was_valid_out\[5\][0] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_3362_ _1795_ _1794_ net1244 _1790_ net1235 VPWR VGND sg13g2_a22oi_1
XFILLER_44_1018 VPWR VGND sg13g2_decap_8
X_5101_ VPWR _0090_ _0798_ VGND sg13g2_inv_1
X_6081_ net198 VGND VPWR _0131_ s0.shift_out\[11\][0] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_3293_ _1731_ VPWR _1732_ VGND _1727_ _1730_ sg13g2_o21ai_1
X_5032_ _0737_ _0736_ net1244 _0732_ net1235 VPWR VGND sg13g2_a22oi_1
X_5934_ _1548_ net1023 _1547_ VPWR VGND sg13g2_nand2b_1
X_5865_ net1013 net1071 _1486_ VPWR VGND sg13g2_nor2b_1
X_4816_ _0540_ VPWR _0541_ VGND net1305 net450 sg13g2_o21ai_1
X_5796_ _1366_ _1421_ net1280 _1422_ VPWR VGND sg13g2_nand3_1
X_4747_ VPWR _0058_ _0476_ VGND sg13g2_inv_1
X_4678_ net924 VPWR _0417_ VGND net321 net1165 sg13g2_o21ai_1
X_3629_ s0.data_out\[4\]\[4\] s0.data_out\[3\]\[4\] net979 _2038_ VPWR VGND sg13g2_mux2_1
XFILLER_0_215 VPWR VGND sg13g2_decap_8
XFILLER_49_709 VPWR VGND sg13g2_decap_8
XFILLER_17_617 VPWR VGND sg13g2_fill_1
XFILLER_29_499 VPWR VGND sg13g2_decap_8
XFILLER_24_160 VPWR VGND sg13g2_fill_2
XFILLER_40_653 VPWR VGND sg13g2_decap_8
XFILLER_9_816 VPWR VGND sg13g2_decap_8
XFILLER_24_193 VPWR VGND sg13g2_fill_1
XFILLER_40_686 VPWR VGND sg13g2_decap_8
XFILLER_40_664 VPWR VGND sg13g2_fill_2
XFILLER_8_304 VPWR VGND sg13g2_fill_1
XFILLER_0_782 VPWR VGND sg13g2_decap_8
XFILLER_48_731 VPWR VGND sg13g2_decap_8
XFILLER_36_959 VPWR VGND sg13g2_decap_8
XFILLER_35_436 VPWR VGND sg13g2_fill_2
XFILLER_35_425 VPWR VGND sg13g2_decap_8
X_3980_ _2353_ net951 _2352_ VPWR VGND sg13g2_nand2b_1
XFILLER_16_683 VPWR VGND sg13g2_fill_2
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
X_5650_ s0.data_out\[10\]\[2\] s0.data_out\[9\]\[2\] net1043 _1295_ VPWR VGND sg13g2_mux2_1
X_4601_ _0344_ VPWR _0345_ VGND _0340_ _0343_ sg13g2_o21ai_1
XFILLER_31_664 VPWR VGND sg13g2_decap_8
XFILLER_31_686 VPWR VGND sg13g2_fill_1
X_5581_ _1235_ VPWR _1236_ VGND net1038 _1229_ sg13g2_o21ai_1
X_4532_ net1262 _2821_ _0285_ VPWR VGND sg13g2_nor2_1
XFILLER_7_40 VPWR VGND sg13g2_fill_2
XFILLER_8_893 VPWR VGND sg13g2_decap_8
X_4463_ VPWR _0031_ _2782_ VGND sg13g2_inv_1
Xhold304 s0.data_new_delayed\[2\] VPWR VGND net600 sg13g2_dlygate4sd3_1
Xhold315 s0.data_out\[2\]\[2\] VPWR VGND net611 sg13g2_dlygate4sd3_1
X_3414_ _1841_ net533 net997 VPWR VGND sg13g2_nand2b_1
X_6202_ net66 VGND VPWR _0252_ s0.data_out\[1\]\[2\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_4394_ VGND VPWR net1183 _2721_ _2722_ _2664_ sg13g2_a21oi_1
X_6133_ net142 VGND VPWR _0183_ s0.data_out\[7\]\[5\] clknet_leaf_16_clk sg13g2_dfrbpq_2
X_3345_ _1778_ net1000 _1777_ VPWR VGND sg13g2_nand2b_1
X_6064_ net216 VGND VPWR _0114_ s0.data_out\[12\]\[3\] clknet_leaf_25_clk sg13g2_dfrbpq_2
X_3276_ _1713_ _1716_ net1324 _1717_ VPWR VGND sg13g2_nand3_1
X_6214__162 VPWR VGND net162 sg13g2_tiehi
XFILLER_39_753 VPWR VGND sg13g2_fill_2
X_5015_ VPWR VGND _0652_ net1282 _0719_ net1277 _0720_ _0716_ sg13g2_a221oi_1
XFILLER_38_285 VPWR VGND sg13g2_decap_8
XFILLER_42_929 VPWR VGND sg13g2_decap_8
XFILLER_26_49 VPWR VGND sg13g2_decap_8
X_5917_ _1531_ VPWR _1532_ VGND _1527_ _1530_ sg13g2_o21ai_1
XFILLER_41_439 VPWR VGND sg13g2_decap_8
XFILLER_35_992 VPWR VGND sg13g2_decap_8
XFILLER_42_48 VPWR VGND sg13g2_decap_8
X_5848_ _1469_ VPWR _1472_ VGND net326 net1021 sg13g2_o21ai_1
X_5779_ VPWR _0160_ net543 VGND sg13g2_inv_1
XFILLER_21_196 VPWR VGND sg13g2_fill_2
XFILLER_5_318 VPWR VGND sg13g2_fill_1
XFILLER_27_1002 VPWR VGND sg13g2_decap_8
XFILLER_49_506 VPWR VGND sg13g2_decap_8
XFILLER_1_557 VPWR VGND sg13g2_decap_8
XFILLER_17_403 VPWR VGND sg13g2_fill_1
XFILLER_17_436 VPWR VGND sg13g2_fill_2
XFILLER_29_285 VPWR VGND sg13g2_decap_8
XFILLER_45_767 VPWR VGND sg13g2_decap_8
XFILLER_17_458 VPWR VGND sg13g2_fill_1
XFILLER_17_469 VPWR VGND sg13g2_fill_1
XFILLER_32_406 VPWR VGND sg13g2_fill_1
XFILLER_44_277 VPWR VGND sg13g2_decap_8
XFILLER_32_428 VPWR VGND sg13g2_fill_1
XFILLER_41_940 VPWR VGND sg13g2_decap_8
XFILLER_34_1028 VPWR VGND sg13g2_fill_1
XFILLER_40_494 VPWR VGND sg13g2_fill_1
XFILLER_8_167 VPWR VGND sg13g2_fill_2
XFILLER_8_156 VPWR VGND sg13g2_decap_8
X_6157__116 VPWR VGND net116 sg13g2_tiehi
XFILLER_5_874 VPWR VGND sg13g2_decap_8
XFILLER_4_340 VPWR VGND sg13g2_decap_8
XFILLER_4_373 VPWR VGND sg13g2_decap_4
X_3130_ net1228 net1010 _1585_ VPWR VGND sg13g2_nor2b_1
XFILLER_36_789 VPWR VGND sg13g2_fill_1
XFILLER_17_970 VPWR VGND sg13g2_decap_8
X_3963_ VGND VPWR _2338_ net590 net1295 sg13g2_or2_1
X_3894_ _2263_ _2278_ _2279_ VPWR VGND sg13g2_nor2b_1
X_5702_ net1069 net1273 net1224 _0145_ VPWR VGND sg13g2_mux2_1
X_5633_ VPWR _0140_ _1280_ VGND sg13g2_inv_1
X_5564_ net1265 _1197_ _1221_ VPWR VGND sg13g2_nor2_1
X_4515_ _2830_ net1170 _2792_ _2831_ VPWR VGND sg13g2_a21o_1
Xhold101 _2304_ VPWR VGND net397 sg13g2_dlygate4sd3_1
Xhold134 s0.data_out\[13\]\[4\] VPWR VGND net430 sg13g2_dlygate4sd3_1
Xhold112 s0.was_valid_out\[12\][0] VPWR VGND net408 sg13g2_dlygate4sd3_1
Xhold123 s0.data_out\[7\]\[1\] VPWR VGND net419 sg13g2_dlygate4sd3_1
X_5495_ VGND VPWR net1081 net429 _1156_ _1155_ sg13g2_a21oi_1
Xhold145 s0.data_out\[3\]\[4\] VPWR VGND net441 sg13g2_dlygate4sd3_1
X_4446_ _2767_ VPWR _2768_ VGND net1287 net475 sg13g2_o21ai_1
Xhold156 s0.data_out\[11\]\[0\] VPWR VGND net452 sg13g2_dlygate4sd3_1
Xhold167 s0.data_out\[5\]\[1\] VPWR VGND net463 sg13g2_dlygate4sd3_1
X_4377_ _2704_ net1179 _2656_ _2705_ VPWR VGND sg13g2_a21o_1
Xhold178 s0.data_out\[15\]\[4\] VPWR VGND net474 sg13g2_dlygate4sd3_1
Xhold189 _1732_ VPWR VGND net485 sg13g2_dlygate4sd3_1
X_3328_ VGND VPWR _1683_ _1761_ _1762_ net1004 sg13g2_a21oi_1
X_6116_ net160 VGND VPWR _0166_ s0.data_out\[8\]\[0\] clknet_leaf_23_clk sg13g2_dfrbpq_2
X_3259_ net1004 VPWR _1702_ VGND net1230 net995 sg13g2_o21ai_1
XFILLER_39_550 VPWR VGND sg13g2_fill_1
X_6047_ net235 VGND VPWR net347 s0.was_valid_out\[13\][0] clknet_leaf_27_clk sg13g2_dfrbpq_2
XFILLER_2_1015 VPWR VGND sg13g2_decap_8
XFILLER_27_767 VPWR VGND sg13g2_decap_8
XFILLER_27_778 VPWR VGND sg13g2_fill_1
XFILLER_14_406 VPWR VGND sg13g2_decap_8
XFILLER_26_277 VPWR VGND sg13g2_fill_1
XFILLER_41_225 VPWR VGND sg13g2_fill_1
XFILLER_10_612 VPWR VGND sg13g2_fill_2
XFILLER_2_833 VPWR VGND sg13g2_decap_8
XFILLER_49_325 VPWR VGND sg13g2_decap_8
XFILLER_45_542 VPWR VGND sg13g2_fill_2
X_6204__40 VPWR VGND net40 sg13g2_tiehi
XFILLER_32_236 VPWR VGND sg13g2_fill_1
XFILLER_13_461 VPWR VGND sg13g2_fill_2
X_5280_ VGND VPWR net1117 _0960_ _0961_ _0910_ sg13g2_a21oi_1
X_4300_ net1178 net1073 _2636_ VPWR VGND sg13g2_nor2b_1
X_6170__102 VPWR VGND net102 sg13g2_tiehi
X_4231_ _2570_ VPWR _2571_ VGND net1198 _2479_ sg13g2_o21ai_1
XFILLER_4_85 VPWR VGND sg13g2_decap_4
X_4162_ _2509_ _2511_ _2512_ VPWR VGND sg13g2_nor2_1
XFILLER_49_870 VPWR VGND sg13g2_decap_8
X_3113_ s0.data_out\[8\]\[5\] s0.data_out\[7\]\[5\] net1021 _1570_ VPWR VGND sg13g2_mux2_1
X_4093_ VPWR _2452_ net1128 VGND sg13g2_inv_1
X_4995_ VGND VPWR _0610_ _0700_ _0701_ net1139 sg13g2_a21oi_1
XFILLER_24_759 VPWR VGND sg13g2_fill_2
X_3946_ net952 VPWR _2323_ VGND _2321_ _2322_ sg13g2_o21ai_1
XFILLER_17_1012 VPWR VGND sg13g2_decap_8
X_3877_ VGND VPWR _2262_ _2259_ net1239 sg13g2_or2_1
XFILLER_20_976 VPWR VGND sg13g2_decap_8
X_5616_ _1265_ VPWR _1266_ VGND net1341 net436 sg13g2_o21ai_1
X_5547_ s0.data_out\[11\]\[6\] s0.data_out\[10\]\[6\] net1085 _1204_ VPWR VGND sg13g2_mux2_1
X_5478_ net1079 net1067 _1141_ VPWR VGND sg13g2_nor2b_1
X_4429_ _2749_ _2752_ net1287 _2753_ VPWR VGND sg13g2_nand3_1
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_47_829 VPWR VGND sg13g2_decap_8
XFILLER_15_715 VPWR VGND sg13g2_decap_8
X_6198__72 VPWR VGND net72 sg13g2_tiehi
X_6008__277 VPWR VGND net277 sg13g2_tiehi
XFILLER_10_431 VPWR VGND sg13g2_decap_8
XFILLER_10_442 VPWR VGND sg13g2_fill_1
XFILLER_22_280 VPWR VGND sg13g2_decap_4
XFILLER_7_936 VPWR VGND sg13g2_decap_8
X_6154__119 VPWR VGND net119 sg13g2_tiehi
XFILLER_37_317 VPWR VGND sg13g2_fill_2
XFILLER_46_873 VPWR VGND sg13g2_decap_8
X_4780_ s0.data_out\[17\]\[4\] s0.data_out\[16\]\[4\] net1151 _0509_ VPWR VGND sg13g2_mux2_1
X_3800_ VGND VPWR _2117_ _2190_ _2191_ net961 sg13g2_a21oi_1
XFILLER_33_556 VPWR VGND sg13g2_fill_2
XFILLER_14_781 VPWR VGND sg13g2_fill_2
XFILLER_20_228 VPWR VGND sg13g2_decap_8
X_3731_ net1284 _2127_ _2128_ VPWR VGND sg13g2_nor2b_1
Xclkload10 VPWR clkload10/Y clknet_leaf_25_clk VGND sg13g2_inv_1
X_3662_ _2066_ VPWR _2067_ VGND net1297 net437 sg13g2_o21ai_1
X_5401_ VGND VPWR net1102 _1069_ _1070_ _1014_ sg13g2_a21oi_1
X_3593_ VGND VPWR net980 _2001_ _2002_ _1959_ sg13g2_a21oi_1
X_5332_ net1088 net1074 _1009_ VPWR VGND sg13g2_nor2b_1
X_6098__180 VPWR VGND net180 sg13g2_tiehi
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_5263_ _0944_ net1108 net504 VPWR VGND sg13g2_nand2_1
X_5194_ net936 VPWR _0885_ VGND s0.was_valid_out\[12\][0] s0.valid_out\[13\][0] sg13g2_o21ai_1
X_4214_ net1195 s0.data_out\[20\]\[6\] _2556_ VPWR VGND sg13g2_and2_1
X_4145_ VGND VPWR net1214 net912 net6 _2499_ sg13g2_a21oi_1
XFILLER_29_829 VPWR VGND sg13g2_decap_8
XFILLER_28_317 VPWR VGND sg13g2_decap_4
XFILLER_28_328 VPWR VGND sg13g2_fill_1
XFILLER_28_339 VPWR VGND sg13g2_decap_8
X_4076_ _2437_ _2474_ _2422_ VPWR VGND sg13g2_nand2b_1
XFILLER_36_372 VPWR VGND sg13g2_decap_8
XFILLER_24_534 VPWR VGND sg13g2_decap_8
XFILLER_11_206 VPWR VGND sg13g2_fill_2
X_4978_ s0.data_out\[14\]\[5\] s0.data_out\[15\]\[5\] net1143 _0686_ VPWR VGND sg13g2_mux2_1
Xclkload4 clknet_leaf_36_clk clkload4/X VPWR VGND sg13g2_buf_8
X_3929_ net942 net1065 _2308_ VPWR VGND sg13g2_nor2b_1
X_6195__75 VPWR VGND net75 sg13g2_tiehi
XFILLER_4_928 VPWR VGND sg13g2_decap_8
Xfanout1228 net1230 net1228 VPWR VGND sg13g2_buf_8
Xfanout1206 net1207 net1206 VPWR VGND sg13g2_buf_8
Xfanout1217 net1218 net1217 VPWR VGND sg13g2_buf_2
Xfanout1239 net1241 net1239 VPWR VGND sg13g2_buf_8
XFILLER_47_626 VPWR VGND sg13g2_decap_8
X_6014__270 VPWR VGND net270 sg13g2_tiehi
XFILLER_15_501 VPWR VGND sg13g2_decap_4
XFILLER_27_372 VPWR VGND sg13g2_fill_1
XFILLER_42_342 VPWR VGND sg13g2_decap_8
XFILLER_15_578 VPWR VGND sg13g2_decap_8
XFILLER_43_898 VPWR VGND sg13g2_decap_8
XFILLER_11_740 VPWR VGND sg13g2_fill_1
XFILLER_7_744 VPWR VGND sg13g2_fill_1
XFILLER_6_221 VPWR VGND sg13g2_fill_1
X_6021__263 VPWR VGND net263 sg13g2_tiehi
XFILLER_6_298 VPWR VGND sg13g2_decap_8
XFILLER_3_950 VPWR VGND sg13g2_decap_8
XFILLER_38_659 VPWR VGND sg13g2_decap_8
Xheichips25_top_sorter_13 VPWR VGND uio_oe[4] sg13g2_tielo
XFILLER_46_670 VPWR VGND sg13g2_decap_8
X_5950_ net221 VGND VPWR _0000_ s0.module0.bubble clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_1_86 VPWR VGND sg13g2_fill_2
XFILLER_19_862 VPWR VGND sg13g2_fill_2
X_4901_ _0618_ _0617_ net1244 _0613_ net1235 VPWR VGND sg13g2_a22oi_1
X_5881_ net1012 s0.data_out\[7\]\[3\] _1500_ VPWR VGND sg13g2_and2_1
X_4832_ _0554_ VPWR _0555_ VGND net1317 net422 sg13g2_o21ai_1
XFILLER_21_526 VPWR VGND sg13g2_decap_8
X_4763_ _0492_ net1161 _0491_ VPWR VGND sg13g2_nand2b_1
X_3714_ net963 net1046 _2112_ VPWR VGND sg13g2_nor2b_1
X_4694_ net1144 net1069 _0430_ VPWR VGND sg13g2_nor2b_1
X_3645_ net1227 net967 _2052_ VPWR VGND sg13g2_nor2b_1
X_6192__78 VPWR VGND net78 sg13g2_tiehi
X_3576_ VGND VPWR _1907_ _1986_ _1987_ net983 sg13g2_a21oi_1
X_5315_ net298 net1209 _0995_ _0107_ VPWR VGND sg13g2_nor3_1
X_5246_ VPWR _0104_ _0929_ VGND sg13g2_inv_1
Xhold16 s0.module0.bubble VPWR VGND net312 sg13g2_dlygate4sd3_1
Xhold38 s0.data_out\[0\]\[7\] VPWR VGND net334 sg13g2_dlygate4sd3_1
Xhold27 s0.was_valid_out\[19\][0] VPWR VGND net323 sg13g2_dlygate4sd3_1
X_5177_ _0870_ net1251 _0865_ VPWR VGND sg13g2_nand2_1
Xhold49 s0.data_out\[0\]\[2\] VPWR VGND net345 sg13g2_dlygate4sd3_1
X_4128_ VPWR _2487_ s0.data_out\[13\]\[2\] VGND sg13g2_inv_1
X_4059_ _2421_ VPWR _2422_ VGND _2465_ net1049 sg13g2_o21ai_1
XFILLER_45_59 VPWR VGND sg13g2_fill_1
XFILLER_25_843 VPWR VGND sg13g2_fill_2
XFILLER_12_504 VPWR VGND sg13g2_decap_8
XFILLER_24_364 VPWR VGND sg13g2_decap_8
XFILLER_24_397 VPWR VGND sg13g2_fill_2
XFILLER_20_570 VPWR VGND sg13g2_fill_1
XFILLER_10_62 VPWR VGND sg13g2_decap_8
Xfanout1003 s0.shift_out\[6\][0] net1003 VPWR VGND sg13g2_buf_1
XFILLER_10_84 VPWR VGND sg13g2_fill_1
XFILLER_48_913 VPWR VGND sg13g2_decap_8
Xfanout1014 s0.shift_out\[7\][0] net1014 VPWR VGND sg13g2_buf_8
Xfanout1025 net1026 net1025 VPWR VGND sg13g2_buf_8
XFILLER_0_964 VPWR VGND sg13g2_decap_8
Xfanout1047 net1048 net1047 VPWR VGND sg13g2_buf_8
Xfanout1036 net1037 net1036 VPWR VGND sg13g2_buf_8
Xfanout1069 net1072 net1069 VPWR VGND sg13g2_buf_8
Xfanout1058 net1060 net1058 VPWR VGND sg13g2_buf_2
XFILLER_47_456 VPWR VGND sg13g2_decap_4
XFILLER_19_71 VPWR VGND sg13g2_decap_4
XFILLER_47_489 VPWR VGND sg13g2_decap_8
XFILLER_15_342 VPWR VGND sg13g2_fill_1
X_6088__190 VPWR VGND net190 sg13g2_tiehi
XFILLER_43_695 VPWR VGND sg13g2_decap_4
XFILLER_30_323 VPWR VGND sg13g2_fill_1
XFILLER_30_389 VPWR VGND sg13g2_fill_2
X_3430_ s0.data_out\[4\]\[4\] s0.data_out\[5\]\[4\] net997 _1855_ VPWR VGND sg13g2_mux2_1
X_3361_ VGND VPWR net1004 _1793_ _1794_ _1755_ sg13g2_a21oi_1
X_5100_ _0797_ VPWR _0798_ VGND net1320 net386 sg13g2_o21ai_1
X_6095__183 VPWR VGND net183 sg13g2_tiehi
X_6080_ net199 VGND VPWR _0130_ s0.data_out\[11\]\[7\] clknet_leaf_20_clk sg13g2_dfrbpq_2
X_5031_ VGND VPWR net1139 _0735_ _0736_ _0694_ sg13g2_a21oi_1
X_3292_ VGND VPWR _1731_ net484 net1324 sg13g2_or2_1
XFILLER_39_979 VPWR VGND sg13g2_decap_8
XFILLER_47_990 VPWR VGND sg13g2_decap_8
XFILLER_25_139 VPWR VGND sg13g2_decap_8
X_5933_ VGND VPWR net1014 _1546_ _1547_ _1501_ sg13g2_a21oi_1
XFILLER_22_824 VPWR VGND sg13g2_fill_1
X_5864_ VGND VPWR _1418_ _1484_ _1485_ net1023 sg13g2_a21oi_1
XFILLER_34_673 VPWR VGND sg13g2_fill_1
XFILLER_34_695 VPWR VGND sg13g2_fill_2
X_4815_ _0536_ _0539_ net1317 _0540_ VPWR VGND sg13g2_nand3_1
X_5795_ _1421_ net1035 _1420_ VPWR VGND sg13g2_nand2b_1
X_4746_ _0475_ VPWR _0476_ VGND net342 _0474_ sg13g2_o21ai_1
X_4677_ net1146 _0412_ _0416_ VPWR VGND sg13g2_nor2_1
X_3628_ _2036_ VPWR _2037_ VGND net1263 _2017_ sg13g2_o21ai_1
XFILLER_1_739 VPWR VGND sg13g2_decap_8
X_3559_ s0.data_out\[3\]\[4\] s0.data_out\[4\]\[4\] net987 _1972_ VPWR VGND sg13g2_mux2_1
XFILLER_48_209 VPWR VGND sg13g2_fill_1
X_5229_ _0914_ VPWR _0915_ VGND _0910_ _0913_ sg13g2_o21ai_1
XFILLER_45_949 VPWR VGND sg13g2_decap_8
XFILLER_44_426 VPWR VGND sg13g2_decap_8
XFILLER_24_172 VPWR VGND sg13g2_decap_4
XFILLER_25_695 VPWR VGND sg13g2_decap_4
XFILLER_12_345 VPWR VGND sg13g2_decap_8
XFILLER_21_50 VPWR VGND sg13g2_fill_1
XFILLER_48_710 VPWR VGND sg13g2_decap_8
XFILLER_0_761 VPWR VGND sg13g2_decap_8
XFILLER_48_787 VPWR VGND sg13g2_decap_8
XFILLER_43_492 VPWR VGND sg13g2_fill_2
X_4600_ VGND VPWR _0344_ net570 net1303 sg13g2_or2_1
XFILLER_30_164 VPWR VGND sg13g2_decap_4
XFILLER_30_197 VPWR VGND sg13g2_fill_2
X_5580_ net934 VPWR _1235_ VGND s0.was_valid_out\[9\][0] net1085 sg13g2_o21ai_1
X_4531_ net1248 _0277_ _0284_ VPWR VGND sg13g2_nor2_1
XFILLER_7_96 VPWR VGND sg13g2_decap_4
Xhold316 s0.data_out\[12\]\[2\] VPWR VGND net612 sg13g2_dlygate4sd3_1
X_4462_ _2781_ VPWR _2782_ VGND net1289 net414 sg13g2_o21ai_1
Xhold305 s0.valid_out\[15\][0] VPWR VGND net601 sg13g2_dlygate4sd3_1
X_3413_ VPWR _0203_ _1840_ VGND sg13g2_inv_1
X_6201_ net68 VGND VPWR _0251_ s0.data_out\[1\]\[1\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_4393_ s0.data_out\[20\]\[4\] s0.data_out\[19\]\[4\] net1188 _2721_ VPWR VGND sg13g2_mux2_1
X_6132_ net143 VGND VPWR _0182_ s0.data_out\[7\]\[4\] clknet_leaf_16_clk sg13g2_dfrbpq_2
X_3344_ VGND VPWR net991 _1776_ _1777_ _1715_ sg13g2_a21oi_1
XFILLER_30_0 VPWR VGND sg13g2_decap_8
X_6063_ net217 VGND VPWR _0113_ s0.data_out\[12\]\[2\] clknet_leaf_27_clk sg13g2_dfrbpq_2
X_3275_ net1000 VPWR _1716_ VGND _1714_ _1715_ sg13g2_o21ai_1
X_5014_ _0719_ net1138 _0718_ VPWR VGND sg13g2_nand2b_1
XFILLER_26_415 VPWR VGND sg13g2_fill_1
XFILLER_42_908 VPWR VGND sg13g2_decap_8
XFILLER_26_448 VPWR VGND sg13g2_decap_8
X_5916_ VGND VPWR _1531_ net595 net1342 sg13g2_or2_1
XFILLER_41_429 VPWR VGND sg13g2_fill_1
XFILLER_35_971 VPWR VGND sg13g2_decap_8
XFILLER_22_643 VPWR VGND sg13g2_decap_8
X_5847_ _1470_ VPWR _1471_ VGND net1029 _1349_ sg13g2_o21ai_1
X_5778_ _1405_ VPWR _1406_ VGND _1401_ _1404_ sg13g2_o21ai_1
XFILLER_10_838 VPWR VGND sg13g2_decap_4
X_4729_ VGND VPWR _0461_ net582 net1306 sg13g2_or2_1
XFILLER_1_536 VPWR VGND sg13g2_decap_8
XFILLER_18_927 VPWR VGND sg13g2_decap_4
XFILLER_45_746 VPWR VGND sg13g2_decap_8
XFILLER_44_256 VPWR VGND sg13g2_decap_8
XFILLER_16_61 VPWR VGND sg13g2_decap_8
XFILLER_13_643 VPWR VGND sg13g2_decap_8
X_6085__193 VPWR VGND net193 sg13g2_tiehi
XFILLER_13_654 VPWR VGND sg13g2_fill_1
XFILLER_41_996 VPWR VGND sg13g2_decap_8
XFILLER_9_636 VPWR VGND sg13g2_fill_1
XFILLER_8_146 VPWR VGND sg13g2_fill_1
XFILLER_32_93 VPWR VGND sg13g2_decap_4
XFILLER_5_853 VPWR VGND sg13g2_decap_8
X_6092__186 VPWR VGND net186 sg13g2_tiehi
XFILLER_48_584 VPWR VGND sg13g2_decap_8
X_5958__59 VPWR VGND net59 sg13g2_tiehi
X_3962_ net1295 VPWR _2337_ VGND net929 _2336_ sg13g2_o21ai_1
X_5701_ net1073 net1281 net1223 _0144_ VPWR VGND sg13g2_mux2_1
X_3893_ _2272_ VPWR _2278_ VGND _2268_ _2274_ sg13g2_o21ai_1
X_5632_ _1279_ VPWR _1280_ VGND net1346 net481 sg13g2_o21ai_1
XFILLER_32_996 VPWR VGND sg13g2_decap_8
X_5563_ net1252 _1217_ _1220_ VPWR VGND sg13g2_nor2_1
X_4514_ s0.data_out\[19\]\[6\] s0.data_out\[18\]\[6\] net1176 _2830_ VPWR VGND sg13g2_mux2_1
Xhold102 s0.was_valid_out\[8\][0] VPWR VGND net398 sg13g2_dlygate4sd3_1
Xhold135 s0.data_out\[15\]\[1\] VPWR VGND net431 sg13g2_dlygate4sd3_1
Xhold113 _0109_ VPWR VGND net409 sg13g2_dlygate4sd3_1
Xhold124 s0.data_out\[3\]\[2\] VPWR VGND net420 sg13g2_dlygate4sd3_1
X_5494_ net1081 net1059 _1155_ VPWR VGND sg13g2_nor2b_1
Xhold157 s0.was_valid_out\[9\][0] VPWR VGND net453 sg13g2_dlygate4sd3_1
Xhold146 s0.data_out\[9\]\[4\] VPWR VGND net442 sg13g2_dlygate4sd3_1
X_4445_ _2763_ _2766_ net1287 _2767_ VPWR VGND sg13g2_nand3_1
Xhold168 s0.data_out\[19\]\[1\] VPWR VGND net464 sg13g2_dlygate4sd3_1
X_4376_ s0.data_out\[20\]\[3\] s0.data_out\[19\]\[3\] net1186 _2704_ VPWR VGND sg13g2_mux2_1
Xhold179 s0.data_out\[19\]\[2\] VPWR VGND net475 sg13g2_dlygate4sd3_1
X_6115_ net161 VGND VPWR _0165_ s0.valid_out\[8\][0] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_3327_ _1761_ s0.data_out\[5\]\[7\] net1009 VPWR VGND sg13g2_nand2b_1
XFILLER_37_49 VPWR VGND sg13g2_fill_1
X_3258_ net1325 net309 _0187_ VPWR VGND sg13g2_and2_1
X_6046_ net236 VGND VPWR _0096_ s0.genblk1\[13\].modules.bubble clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
X_3189_ _1636_ s0.data_out\[6\]\[6\] net1020 VPWR VGND sg13g2_nand2b_1
XFILLER_27_724 VPWR VGND sg13g2_fill_2
XFILLER_14_429 VPWR VGND sg13g2_decap_4
XFILLER_35_790 VPWR VGND sg13g2_decap_4
XFILLER_23_985 VPWR VGND sg13g2_decap_8
XFILLER_2_812 VPWR VGND sg13g2_decap_8
XFILLER_49_304 VPWR VGND sg13g2_decap_8
XFILLER_2_889 VPWR VGND sg13g2_decap_8
XFILLER_49_348 VPWR VGND sg13g2_fill_2
XFILLER_49_359 VPWR VGND sg13g2_decap_8
XFILLER_40_1022 VPWR VGND sg13g2_decap_8
XFILLER_27_82 VPWR VGND sg13g2_fill_2
XFILLER_41_782 VPWR VGND sg13g2_decap_4
XFILLER_14_996 VPWR VGND sg13g2_decap_8
XFILLER_9_466 VPWR VGND sg13g2_decap_8
X_4230_ _2570_ net1198 net490 VPWR VGND sg13g2_nand2_1
XFILLER_4_20 VPWR VGND sg13g2_fill_2
X_4161_ _2510_ VPWR _2511_ VGND net1195 _2503_ sg13g2_o21ai_1
X_3112_ _1569_ net1020 net589 VPWR VGND sg13g2_nand2_1
X_4092_ VPWR _2451_ net1105 VGND sg13g2_inv_1
XFILLER_36_532 VPWR VGND sg13g2_decap_8
X_4994_ _0700_ s0.data_out\[14\]\[7\] net1142 VPWR VGND sg13g2_nand2b_1
X_3945_ net942 net1057 _2322_ VPWR VGND sg13g2_nor2b_1
X_3876_ VGND VPWR _2261_ _2255_ net1232 sg13g2_or2_1
XFILLER_20_966 VPWR VGND sg13g2_fill_1
X_5615_ _1261_ _1264_ net1341 _1265_ VPWR VGND sg13g2_nand3_1
X_5546_ _1203_ net1086 net521 VPWR VGND sg13g2_nand2_1
X_5477_ VGND VPWR _1062_ _1139_ _1140_ net1090 sg13g2_a21oi_1
X_4428_ net1181 VPWR _2752_ VGND _2750_ _2751_ sg13g2_o21ai_1
X_4359_ _2687_ VPWR _2688_ VGND _2683_ _2686_ sg13g2_o21ai_1
XFILLER_47_808 VPWR VGND sg13g2_decap_8
XFILLER_24_1028 VPWR VGND sg13g2_fill_1
X_6029_ net254 VGND VPWR _0079_ s0.data_out\[15\]\[4\] clknet_leaf_23_clk sg13g2_dfrbpq_2
XFILLER_27_543 VPWR VGND sg13g2_decap_4
X_6147__127 VPWR VGND net127 sg13g2_tiehi
XFILLER_42_502 VPWR VGND sg13g2_fill_2
XFILLER_42_524 VPWR VGND sg13g2_decap_8
XFILLER_14_226 VPWR VGND sg13g2_fill_1
XFILLER_7_915 VPWR VGND sg13g2_decap_8
XFILLER_22_292 VPWR VGND sg13g2_fill_2
XFILLER_11_988 VPWR VGND sg13g2_decap_8
XFILLER_6_447 VPWR VGND sg13g2_fill_2
XFILLER_2_675 VPWR VGND sg13g2_decap_8
XFILLER_49_112 VPWR VGND sg13g2_decap_8
XFILLER_49_134 VPWR VGND sg13g2_decap_8
XFILLER_49_189 VPWR VGND sg13g2_decap_8
XFILLER_49_167 VPWR VGND sg13g2_decap_8
Xfanout990 net993 net990 VPWR VGND sg13g2_buf_8
XFILLER_46_852 VPWR VGND sg13g2_decap_8
XFILLER_38_92 VPWR VGND sg13g2_decap_8
XFILLER_45_373 VPWR VGND sg13g2_fill_1
X_3730_ _2062_ VPWR _2127_ VGND net932 _2126_ sg13g2_o21ai_1
X_3661_ _2062_ _2065_ net1307 _2066_ VPWR VGND sg13g2_nand3_1
Xclkload11 clkload11/Y clknet_leaf_28_clk VPWR VGND sg13g2_inv_8
X_5400_ _1068_ net1088 _1015_ _1069_ VPWR VGND sg13g2_a21o_1
X_3592_ _2000_ net969 _1960_ _2001_ VPWR VGND sg13g2_a21o_1
X_5331_ net1088 s0.data_out\[11\]\[0\] _1008_ VPWR VGND sg13g2_and2_1
X_5262_ VPWR _0106_ net585 VGND sg13g2_inv_1
X_5193_ net1107 _0878_ _0884_ VPWR VGND sg13g2_nor2_1
X_4213_ _0008_ _2551_ _2555_ _2475_ net1217 VPWR VGND sg13g2_a22oi_1
X_4144_ s0.data_out\[21\]\[4\] net912 _2499_ VPWR VGND sg13g2_nor2_1
XFILLER_29_808 VPWR VGND sg13g2_decap_4
X_4075_ _2436_ _2426_ _2435_ _2422_ net1241 VPWR VGND sg13g2_a22oi_1
XFILLER_37_863 VPWR VGND sg13g2_fill_2
XFILLER_34_17 VPWR VGND sg13g2_decap_8
X_4977_ VPWR _0079_ _0685_ VGND sg13g2_inv_1
Xclkload5 clkload5/Y clknet_leaf_37_clk VPWR VGND sg13g2_inv_2
X_3928_ net940 s0.data_out\[0\]\[2\] _2307_ VPWR VGND sg13g2_and2_1
XFILLER_32_590 VPWR VGND sg13g2_fill_1
X_3859_ _2235_ VPWR _2244_ VGND net1273 _2239_ sg13g2_o21ai_1
XFILLER_4_907 VPWR VGND sg13g2_decap_8
XFILLER_3_417 VPWR VGND sg13g2_decap_4
X_5529_ s0.data_out\[11\]\[1\] s0.data_out\[10\]\[1\] net1084 _1186_ VPWR VGND sg13g2_mux2_1
X_6153__120 VPWR VGND net120 sg13g2_tiehi
Xfanout1229 net1230 net1229 VPWR VGND sg13g2_buf_8
Xfanout1218 net1219 net1218 VPWR VGND sg13g2_buf_8
Xfanout1207 s0.valid_out\[21\][0] net1207 VPWR VGND sg13g2_buf_8
XFILLER_46_148 VPWR VGND sg13g2_fill_1
XFILLER_43_877 VPWR VGND sg13g2_decap_8
XFILLER_15_557 VPWR VGND sg13g2_fill_2
X_6160__113 VPWR VGND net113 sg13g2_tiehi
XFILLER_30_505 VPWR VGND sg13g2_decap_8
XFILLER_24_83 VPWR VGND sg13g2_decap_4
XFILLER_10_273 VPWR VGND sg13g2_fill_2
XFILLER_34_7 VPWR VGND sg13g2_decap_8
XFILLER_49_91 VPWR VGND sg13g2_decap_8
XFILLER_49_80 VPWR VGND sg13g2_fill_2
XFILLER_37_104 VPWR VGND sg13g2_fill_1
XFILLER_37_137 VPWR VGND sg13g2_decap_8
Xheichips25_top_sorter_14 VPWR VGND uio_oe[6] sg13g2_tielo
XFILLER_18_340 VPWR VGND sg13g2_fill_1
XFILLER_19_885 VPWR VGND sg13g2_fill_2
X_4900_ VGND VPWR net1148 _0616_ _0617_ _0578_ sg13g2_a21oi_1
X_5880_ _1499_ net918 _1498_ VPWR VGND sg13g2_nand2_1
XFILLER_34_822 VPWR VGND sg13g2_fill_1
X_4831_ _0550_ _0553_ net1317 _0554_ VPWR VGND sg13g2_nand3_1
X_4762_ VGND VPWR net1147 _0490_ _0491_ _0445_ sg13g2_a21oi_1
XFILLER_21_549 VPWR VGND sg13g2_fill_2
X_3713_ VGND VPWR _2020_ _2110_ _2111_ net973 sg13g2_a21oi_1
X_4693_ VGND VPWR _0365_ _0428_ _0429_ net1162 sg13g2_a21oi_1
X_3644_ net973 VPWR _2051_ VGND net1227 net963 sg13g2_o21ai_1
X_3575_ _1986_ s0.data_out\[3\]\[6\] net988 VPWR VGND sg13g2_nand2b_1
X_5314_ VPWR VGND _0977_ _0994_ _0993_ _0964_ _0995_ _0992_ sg13g2_a221oi_1
X_5245_ _0928_ VPWR _0929_ VGND _0924_ _0927_ sg13g2_o21ai_1
Xhold17 s0.genblk1\[7\].modules.bubble VPWR VGND net313 sg13g2_dlygate4sd3_1
Xhold28 _0025_ VPWR VGND net324 sg13g2_dlygate4sd3_1
X_5176_ _0868_ VPWR _0869_ VGND net1265 _0844_ sg13g2_o21ai_1
Xhold39 s0.shift_out\[14\][0] VPWR VGND net335 sg13g2_dlygate4sd3_1
XFILLER_29_638 VPWR VGND sg13g2_decap_8
X_4127_ VPWR _2486_ net386 VGND sg13g2_inv_1
XFILLER_28_126 VPWR VGND sg13g2_fill_1
XFILLER_28_148 VPWR VGND sg13g2_fill_2
XFILLER_43_107 VPWR VGND sg13g2_decap_8
X_4058_ net351 net947 net944 _2421_ VPWR VGND sg13g2_a21o_1
XFILLER_36_192 VPWR VGND sg13g2_fill_1
XFILLER_24_321 VPWR VGND sg13g2_decap_8
XFILLER_20_582 VPWR VGND sg13g2_fill_1
XFILLER_3_247 VPWR VGND sg13g2_fill_1
Xfanout1004 net1007 net1004 VPWR VGND sg13g2_buf_8
Xfanout1015 net1018 net1015 VPWR VGND sg13g2_buf_8
Xfanout1026 s0.shift_out\[8\][0] net1026 VPWR VGND sg13g2_buf_8
Xfanout1037 net343 net1037 VPWR VGND sg13g2_buf_8
XFILLER_0_943 VPWR VGND sg13g2_decap_8
Xfanout1059 net1060 net1059 VPWR VGND sg13g2_buf_8
Xfanout1048 net593 net1048 VPWR VGND sg13g2_buf_8
XFILLER_48_969 VPWR VGND sg13g2_decap_8
XFILLER_19_50 VPWR VGND sg13g2_fill_2
XFILLER_15_310 VPWR VGND sg13g2_fill_2
XFILLER_16_844 VPWR VGND sg13g2_decap_4
XFILLER_31_803 VPWR VGND sg13g2_decap_8
XFILLER_37_1027 VPWR VGND sg13g2_fill_2
XFILLER_35_71 VPWR VGND sg13g2_decap_4
XFILLER_7_531 VPWR VGND sg13g2_fill_2
XFILLER_7_564 VPWR VGND sg13g2_fill_1
X_3360_ _1792_ net995 _1756_ _1793_ VPWR VGND sg13g2_a21o_1
X_5030_ _0734_ net1125 _0695_ _0735_ VPWR VGND sg13g2_a21o_1
X_3291_ net1326 VPWR _1730_ VGND net916 _1729_ sg13g2_o21ai_1
XFILLER_39_958 VPWR VGND sg13g2_decap_8
XFILLER_38_468 VPWR VGND sg13g2_decap_4
XFILLER_19_693 VPWR VGND sg13g2_decap_4
X_5932_ s0.data_out\[8\]\[3\] s0.data_out\[7\]\[3\] net1022 _1546_ VPWR VGND sg13g2_mux2_1
X_5863_ _1484_ net419 net1031 VPWR VGND sg13g2_nand2b_1
X_4814_ net1149 VPWR _0539_ VGND _0537_ _0538_ sg13g2_o21ai_1
X_5794_ VGND VPWR net1030 _1419_ _1420_ _1368_ sg13g2_a21oi_1
XFILLER_33_195 VPWR VGND sg13g2_decap_8
X_4745_ VGND VPWR _0475_ net341 net1305 sg13g2_or2_1
X_4676_ _0413_ VPWR _0415_ VGND net321 net1151 sg13g2_o21ai_1
X_3627_ _1980_ _2035_ net1249 _2036_ VPWR VGND sg13g2_nand3_1
X_6004__281 VPWR VGND net281 sg13g2_tiehi
XFILLER_1_718 VPWR VGND sg13g2_decap_8
X_3558_ VPWR _0217_ _1971_ VGND sg13g2_inv_1
XFILLER_0_206 VPWR VGND sg13g2_fill_2
X_3489_ VGND VPWR net996 _1909_ _1910_ _1870_ sg13g2_a21oi_1
XFILLER_0_239 VPWR VGND sg13g2_decap_8
X_5228_ VGND VPWR _0914_ net507 net1332 sg13g2_or2_1
XFILLER_5_1014 VPWR VGND sg13g2_decap_8
XFILLER_29_402 VPWR VGND sg13g2_fill_2
X_5159_ _0851_ net1114 _0815_ _0852_ VPWR VGND sg13g2_a21o_1
XFILLER_29_435 VPWR VGND sg13g2_decap_8
XFILLER_45_928 VPWR VGND sg13g2_decap_8
XFILLER_44_449 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_36_clk clknet_3_0__leaf_clk clknet_leaf_36_clk VPWR VGND sg13g2_buf_8
X_6011__274 VPWR VGND net274 sg13g2_tiehi
XFILLER_24_162 VPWR VGND sg13g2_fill_1
XFILLER_9_807 VPWR VGND sg13g2_decap_4
XFILLER_0_740 VPWR VGND sg13g2_decap_8
XFILLER_48_766 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_27_clk clknet_3_5__leaf_clk clknet_leaf_27_clk VPWR VGND sg13g2_buf_8
XFILLER_44_983 VPWR VGND sg13g2_decap_8
XFILLER_31_611 VPWR VGND sg13g2_fill_2
XFILLER_31_633 VPWR VGND sg13g2_fill_2
XFILLER_30_132 VPWR VGND sg13g2_decap_4
XFILLER_31_655 VPWR VGND sg13g2_decap_4
X_4530_ VGND VPWR _2777_ _0281_ _0283_ net1254 sg13g2_a21oi_1
X_4461_ _2777_ _2780_ net1289 _2781_ VPWR VGND sg13g2_nand3_1
Xhold306 s0.data_new_delayed\[4\] VPWR VGND net602 sg13g2_dlygate4sd3_1
Xhold317 s0.data_out\[11\]\[3\] VPWR VGND net613 sg13g2_dlygate4sd3_1
X_3412_ _1839_ VPWR _1840_ VGND net1311 net463 sg13g2_o21ai_1
X_6200_ net69 VGND VPWR _0250_ s0.data_out\[1\]\[0\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_4392_ _2720_ _2717_ _2718_ _2719_ VPWR VGND sg13g2_and3_1
X_6131_ net144 VGND VPWR _0181_ s0.data_out\[7\]\[3\] clknet_leaf_15_clk sg13g2_dfrbpq_2
X_3343_ s0.data_out\[6\]\[0\] s0.data_out\[5\]\[0\] net997 _1776_ VPWR VGND sg13g2_mux2_1
X_6062_ net218 VGND VPWR _0112_ s0.data_out\[12\]\[1\] clknet_leaf_25_clk sg13g2_dfrbpq_2
XFILLER_23_0 VPWR VGND sg13g2_fill_1
X_3274_ net991 net1074 _1715_ VPWR VGND sg13g2_nor2b_1
X_5013_ VGND VPWR net1122 _0717_ _0718_ _0654_ sg13g2_a21oi_1
XFILLER_26_29 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_18_clk clknet_3_7__leaf_clk clknet_leaf_18_clk VPWR VGND sg13g2_buf_8
XFILLER_35_950 VPWR VGND sg13g2_decap_8
X_5915_ net1330 VPWR _1530_ VGND net918 _1529_ sg13g2_o21ai_1
XFILLER_41_408 VPWR VGND sg13g2_fill_2
X_5846_ VPWR _1470_ _1469_ VGND sg13g2_inv_1
XFILLER_22_622 VPWR VGND sg13g2_decap_8
XFILLER_21_132 VPWR VGND sg13g2_decap_8
X_5777_ VGND VPWR _1405_ net542 net1342 sg13g2_or2_1
X_4728_ net1306 VPWR _0460_ VGND _2462_ _0459_ sg13g2_o21ai_1
X_4659_ VGND VPWR net1158 _0399_ _0400_ _0335_ sg13g2_a21oi_1
XFILLER_45_725 VPWR VGND sg13g2_decap_8
XFILLER_26_950 VPWR VGND sg13g2_fill_1
XFILLER_33_909 VPWR VGND sg13g2_decap_8
X_5967__49 VPWR VGND net49 sg13g2_tiehi
XFILLER_26_961 VPWR VGND sg13g2_fill_2
XFILLER_26_994 VPWR VGND sg13g2_decap_8
XFILLER_32_419 VPWR VGND sg13g2_decap_8
XFILLER_41_975 VPWR VGND sg13g2_decap_8
XFILLER_9_604 VPWR VGND sg13g2_decap_4
XFILLER_34_1019 VPWR VGND sg13g2_decap_8
XFILLER_40_485 VPWR VGND sg13g2_decap_4
XFILLER_8_136 VPWR VGND sg13g2_fill_2
XFILLER_5_832 VPWR VGND sg13g2_decap_8
XFILLER_48_563 VPWR VGND sg13g2_decap_8
XFILLER_48_541 VPWR VGND sg13g2_fill_2
X_3961_ VGND VPWR net943 net351 _2336_ _2335_ sg13g2_a21oi_1
XFILLER_32_920 VPWR VGND sg13g2_decap_8
XFILLER_32_931 VPWR VGND sg13g2_decap_4
X_5700_ VGND VPWR _1341_ _1343_ _0143_ _1344_ sg13g2_a21oi_1
X_3892_ _2264_ _2272_ _2251_ _2277_ VPWR VGND _2276_ sg13g2_nand4_1
XFILLER_32_975 VPWR VGND sg13g2_decap_8
X_5631_ _1275_ _1278_ net1346 _1279_ VPWR VGND sg13g2_nand3_1
X_5562_ net1256 _1213_ _1219_ VPWR VGND sg13g2_nor2_1
X_4513_ _2829_ net1176 net558 VPWR VGND sg13g2_nand2_1
Xhold103 _0164_ VPWR VGND net399 sg13g2_dlygate4sd3_1
Xhold114 s0.data_out\[19\]\[0\] VPWR VGND net410 sg13g2_dlygate4sd3_1
Xhold125 s0.data_out\[3\]\[1\] VPWR VGND net421 sg13g2_dlygate4sd3_1
X_5493_ VGND VPWR _1095_ _1153_ _1154_ net1093 sg13g2_a21oi_1
X_4444_ net1181 VPWR _2766_ VGND _2764_ _2765_ sg13g2_o21ai_1
Xhold136 s0.data_out\[5\]\[0\] VPWR VGND net432 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_3_2__leaf_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
Xhold158 s0.data_out\[6\]\[3\] VPWR VGND net454 sg13g2_dlygate4sd3_1
Xhold147 s0.data_out\[4\]\[4\] VPWR VGND net443 sg13g2_dlygate4sd3_1
Xhold169 s0.was_valid_out\[6\][0] VPWR VGND net465 sg13g2_dlygate4sd3_1
X_4375_ _2703_ net1186 net567 VPWR VGND sg13g2_nand2_1
X_6001__284 VPWR VGND net284 sg13g2_tiehi
X_3326_ VPWR _0196_ _1760_ VGND sg13g2_inv_1
X_6114_ net163 VGND VPWR net399 s0.was_valid_out\[8\][0] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_6045_ net237 VGND VPWR _0095_ s0.shift_out\[14\][0] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_3257_ _1700_ _1701_ _0186_ VPWR VGND sg13g2_and2_1
XFILLER_27_703 VPWR VGND sg13g2_decap_8
X_3188_ VPWR _0183_ _1635_ VGND sg13g2_inv_1
XFILLER_26_202 VPWR VGND sg13g2_fill_2
XFILLER_22_452 VPWR VGND sg13g2_decap_8
XFILLER_23_964 VPWR VGND sg13g2_decap_8
X_5957__60 VPWR VGND net60 sg13g2_tiehi
XFILLER_34_290 VPWR VGND sg13g2_decap_8
X_5829_ s0.data_out\[9\]\[4\] s0.data_out\[8\]\[4\] net1033 _1455_ VPWR VGND sg13g2_mux2_1
XFILLER_10_625 VPWR VGND sg13g2_decap_8
XFILLER_22_485 VPWR VGND sg13g2_decap_4
XFILLER_2_868 VPWR VGND sg13g2_decap_8
XFILLER_40_1001 VPWR VGND sg13g2_decap_8
XFILLER_45_544 VPWR VGND sg13g2_fill_1
XFILLER_17_246 VPWR VGND sg13g2_decap_8
XFILLER_27_61 VPWR VGND sg13g2_fill_1
XFILLER_27_94 VPWR VGND sg13g2_fill_2
XFILLER_13_452 VPWR VGND sg13g2_decap_4
XFILLER_14_975 VPWR VGND sg13g2_decap_8
XFILLER_25_290 VPWR VGND sg13g2_decap_8
XFILLER_9_434 VPWR VGND sg13g2_decap_8
X_4160_ _2457_ VPWR _2510_ VGND s0.was_valid_out\[20\][0] net1207 sg13g2_o21ai_1
X_3111_ _1506_ _1567_ net1256 _1568_ VPWR VGND sg13g2_nand3_1
X_4091_ net1337 _2450_ VPWR VGND sg13g2_inv_4
XFILLER_48_393 VPWR VGND sg13g2_decap_4
XFILLER_48_382 VPWR VGND sg13g2_fill_2
X_4993_ VPWR _0081_ net563 VGND sg13g2_inv_1
X_3944_ net945 s0.data_out\[0\]\[4\] _2321_ VPWR VGND sg13g2_and2_1
X_3875_ _2260_ _2259_ net1239 _2255_ net1232 VPWR VGND sg13g2_a22oi_1
XFILLER_20_912 VPWR VGND sg13g2_fill_2
XFILLER_31_271 VPWR VGND sg13g2_decap_8
X_5954__63 VPWR VGND net63 sg13g2_tiehi
X_5614_ net1079 VPWR _1264_ VGND _1262_ _1263_ sg13g2_o21ai_1
X_5545_ VGND VPWR net1094 _1201_ _1202_ _1175_ sg13g2_a21oi_1
X_5476_ _1139_ net506 net1096 VPWR VGND sg13g2_nand2b_1
X_4427_ net1167 net1073 _2751_ VPWR VGND sg13g2_nor2b_1
X_4358_ VGND VPWR _2687_ net523 net1288 sg13g2_or2_1
XFILLER_24_1007 VPWR VGND sg13g2_decap_8
X_4289_ net323 net1188 _2627_ VPWR VGND sg13g2_nor2_1
X_3309_ _1745_ VPWR _1746_ VGND net1324 net423 sg13g2_o21ai_1
X_6028_ net255 VGND VPWR _0078_ s0.data_out\[15\]\[3\] clknet_leaf_30_clk sg13g2_dfrbpq_2
XFILLER_27_511 VPWR VGND sg13g2_fill_1
XFILLER_42_536 VPWR VGND sg13g2_decap_8
XFILLER_27_599 VPWR VGND sg13g2_decap_8
XFILLER_42_569 VPWR VGND sg13g2_decap_4
X_6082__197 VPWR VGND net197 sg13g2_tiehi
XFILLER_11_967 VPWR VGND sg13g2_decap_8
XFILLER_2_654 VPWR VGND sg13g2_decap_8
XFILLER_2_643 VPWR VGND sg13g2_decap_4
XFILLER_1_197 VPWR VGND sg13g2_decap_4
XFILLER_38_60 VPWR VGND sg13g2_decap_8
Xfanout991 net992 net991 VPWR VGND sg13g2_buf_2
Xfanout980 net986 net980 VPWR VGND sg13g2_buf_8
XFILLER_46_831 VPWR VGND sg13g2_decap_8
XFILLER_18_544 VPWR VGND sg13g2_fill_2
XFILLER_45_352 VPWR VGND sg13g2_decap_8
XFILLER_45_396 VPWR VGND sg13g2_fill_1
XFILLER_14_783 VPWR VGND sg13g2_fill_1
X_3660_ net971 VPWR _2065_ VGND _2063_ _2064_ sg13g2_o21ai_1
Xclkload12 clkload12/Y clknet_leaf_5_clk VPWR VGND sg13g2_inv_2
X_3591_ s0.data_out\[4\]\[2\] s0.data_out\[3\]\[2\] net979 _2000_ VPWR VGND sg13g2_mux2_1
XFILLER_6_982 VPWR VGND sg13g2_decap_8
X_5330_ _1007_ net938 _1006_ VPWR VGND sg13g2_nand2_1
XFILLER_47_1018 VPWR VGND sg13g2_decap_8
X_5261_ _0942_ VPWR _0943_ VGND _0938_ _0941_ sg13g2_o21ai_1
XFILLER_5_481 VPWR VGND sg13g2_decap_8
X_4212_ net1217 _2554_ _2555_ VPWR VGND sg13g2_nor2_1
X_5192_ _0880_ VPWR _0883_ VGND s0.was_valid_out\[12\][0] net1111 sg13g2_o21ai_1
X_4143_ _2498_ VPWR net5 VGND _2478_ net913 sg13g2_o21ai_1
XFILLER_18_19 VPWR VGND sg13g2_decap_8
X_4074_ _2427_ VPWR _2435_ VGND _2432_ _2434_ sg13g2_o21ai_1
XFILLER_36_396 VPWR VGND sg13g2_fill_2
X_4976_ _0684_ VPWR _0685_ VGND net1322 net474 sg13g2_o21ai_1
XFILLER_20_742 VPWR VGND sg13g2_decap_4
X_3927_ _2306_ net928 _2305_ VPWR VGND sg13g2_nand2_1
Xclkload6 clkload6/Y clknet_leaf_35_clk VPWR VGND sg13g2_inv_2
X_3858_ VPWR VGND _2177_ net1281 _2242_ net1273 _2243_ _2239_ sg13g2_a221oi_1
X_3789_ _2181_ VPWR _2182_ VGND net1300 net424 sg13g2_o21ai_1
X_5528_ net1270 _1184_ _1185_ VPWR VGND sg13g2_nor2_1
X_5459_ net1221 _1119_ _0122_ VPWR VGND sg13g2_nor2_1
Xfanout1219 _2450_ net1219 VPWR VGND sg13g2_buf_8
Xfanout1208 net1210 net1208 VPWR VGND sg13g2_buf_8
XFILLER_47_606 VPWR VGND sg13g2_fill_2
XFILLER_46_105 VPWR VGND sg13g2_fill_2
XFILLER_43_856 VPWR VGND sg13g2_decap_8
XFILLER_24_73 VPWR VGND sg13g2_fill_2
XFILLER_6_234 VPWR VGND sg13g2_fill_2
XFILLER_3_985 VPWR VGND sg13g2_decap_8
XFILLER_1_11 VPWR VGND sg13g2_decap_8
XFILLER_1_44 VPWR VGND sg13g2_fill_2
XFILLER_19_864 VPWR VGND sg13g2_fill_1
Xheichips25_top_sorter_15 VPWR VGND uio_oe[7] sg13g2_tielo
X_4830_ net1149 VPWR _0553_ VGND _0551_ _0552_ sg13g2_o21ai_1
XFILLER_33_388 VPWR VGND sg13g2_decap_4
X_4761_ s0.data_out\[17\]\[3\] s0.data_out\[16\]\[3\] net1151 _0490_ VPWR VGND sg13g2_mux2_1
X_3712_ _2110_ s0.data_out\[2\]\[7\] net977 VPWR VGND sg13g2_nand2b_1
X_4692_ _0428_ net476 net1164 VPWR VGND sg13g2_nand2b_1
XFILLER_14_1017 VPWR VGND sg13g2_decap_8
XFILLER_14_1028 VPWR VGND sg13g2_fill_1
X_3643_ net1309 net311 _0223_ VPWR VGND sg13g2_and2_1
X_3574_ VPWR _0219_ _1985_ VGND sg13g2_inv_1
XFILLER_6_790 VPWR VGND sg13g2_fill_1
X_5313_ _0882_ VPWR _0994_ VGND _0973_ _0975_ sg13g2_o21ai_1
X_6137__138 VPWR VGND net138 sg13g2_tiehi
X_5244_ VGND VPWR _0928_ net599 net1338 sg13g2_or2_1
Xhold18 s0.genblk1\[9\].modules.bubble VPWR VGND net314 sg13g2_dlygate4sd3_1
X_5175_ VGND VPWR _0868_ _0860_ net1256 sg13g2_or2_1
Xhold29 s0.data_out\[18\]\[4\] VPWR VGND net325 sg13g2_dlygate4sd3_1
X_4126_ _2485_ net550 VPWR VGND sg13g2_inv_2
XFILLER_45_17 VPWR VGND sg13g2_decap_4
X_4057_ net1294 net351 _2420_ VPWR VGND sg13g2_nor2_1
XFILLER_37_672 VPWR VGND sg13g2_fill_1
XFILLER_36_171 VPWR VGND sg13g2_decap_4
XFILLER_36_160 VPWR VGND sg13g2_fill_1
XFILLER_25_845 VPWR VGND sg13g2_fill_1
X_4959_ _0666_ _0669_ net1320 _0670_ VPWR VGND sg13g2_nand3_1
XFILLER_24_399 VPWR VGND sg13g2_fill_1
XFILLER_4_749 VPWR VGND sg13g2_decap_4
XFILLER_0_922 VPWR VGND sg13g2_decap_8
Xfanout1016 net1018 net1016 VPWR VGND sg13g2_buf_8
Xfanout1005 net1007 net1005 VPWR VGND sg13g2_buf_8
Xfanout1027 net1029 net1027 VPWR VGND sg13g2_buf_8
Xfanout1038 net1040 net1038 VPWR VGND sg13g2_buf_8
XFILLER_47_414 VPWR VGND sg13g2_decap_8
XFILLER_0_999 VPWR VGND sg13g2_decap_8
Xfanout1049 net1052 net1049 VPWR VGND sg13g2_buf_8
XFILLER_48_948 VPWR VGND sg13g2_decap_8
XFILLER_19_138 VPWR VGND sg13g2_decap_4
XFILLER_43_653 VPWR VGND sg13g2_decap_8
XFILLER_37_1006 VPWR VGND sg13g2_decap_8
XFILLER_30_303 VPWR VGND sg13g2_fill_1
XFILLER_30_314 VPWR VGND sg13g2_fill_2
XFILLER_7_554 VPWR VGND sg13g2_fill_1
XFILLER_3_782 VPWR VGND sg13g2_decap_8
X_3290_ VGND VPWR net991 s0.data_out\[5\]\[2\] _1729_ _1728_ sg13g2_a21oi_1
XFILLER_39_937 VPWR VGND sg13g2_decap_8
XFILLER_38_403 VPWR VGND sg13g2_fill_2
XFILLER_25_4 VPWR VGND sg13g2_decap_8
XFILLER_19_650 VPWR VGND sg13g2_decap_4
XFILLER_18_160 VPWR VGND sg13g2_decap_8
X_5931_ _1545_ net1019 net503 VPWR VGND sg13g2_nand2_1
XFILLER_18_182 VPWR VGND sg13g2_fill_1
XFILLER_18_171 VPWR VGND sg13g2_fill_2
XFILLER_34_653 VPWR VGND sg13g2_decap_4
XFILLER_22_815 VPWR VGND sg13g2_decap_8
X_5862_ VPWR _0166_ _1483_ VGND sg13g2_inv_1
X_4813_ net1134 net1074 _0538_ VPWR VGND sg13g2_nor2b_1
X_5793_ s0.data_out\[9\]\[1\] s0.data_out\[8\]\[1\] net1034 _1419_ VPWR VGND sg13g2_mux2_1
X_6143__131 VPWR VGND net131 sg13g2_tiehi
X_4744_ net1304 VPWR _0474_ VGND net924 _0473_ sg13g2_o21ai_1
X_4675_ VPWR _0414_ _0413_ VGND sg13g2_inv_1
X_3626_ _2035_ net983 _2034_ VPWR VGND sg13g2_nand2b_1
X_3557_ _1970_ VPWR _1971_ VGND net1312 net403 sg13g2_o21ai_1
X_3488_ _1908_ net984 _1871_ _1909_ VPWR VGND sg13g2_a21o_1
X_5227_ net1332 VPWR _0913_ VGND net935 _0912_ sg13g2_o21ai_1
XFILLER_0_229 VPWR VGND sg13g2_fill_2
X_6150__124 VPWR VGND net124 sg13g2_tiehi
X_5158_ s0.data_out\[14\]\[6\] s0.data_out\[13\]\[6\] net1120 _0851_ VPWR VGND sg13g2_mux2_1
XFILLER_45_907 VPWR VGND sg13g2_decap_8
X_5089_ VGND VPWR net1112 net477 _0788_ _0787_ sg13g2_a21oi_1
X_4109_ _2468_ net1012 VPWR VGND sg13g2_inv_2
X_5979__36 VPWR VGND net36 sg13g2_tiehi
XFILLER_16_108 VPWR VGND sg13g2_fill_1
XFILLER_12_303 VPWR VGND sg13g2_fill_2
XFILLER_21_85 VPWR VGND sg13g2_fill_2
XFILLER_43_1010 VPWR VGND sg13g2_decap_8
XFILLER_48_745 VPWR VGND sg13g2_decap_8
XFILLER_47_222 VPWR VGND sg13g2_fill_2
XFILLER_0_796 VPWR VGND sg13g2_decap_8
XFILLER_47_255 VPWR VGND sg13g2_fill_2
XFILLER_36_907 VPWR VGND sg13g2_fill_1
XFILLER_29_981 VPWR VGND sg13g2_decap_8
XFILLER_44_962 VPWR VGND sg13g2_decap_8
X_6127__148 VPWR VGND net148 sg13g2_tiehi
XFILLER_30_188 VPWR VGND sg13g2_fill_2
XFILLER_7_54 VPWR VGND sg13g2_decap_4
XFILLER_11_1009 VPWR VGND sg13g2_decap_8
X_4460_ net1183 VPWR _2780_ VGND _2778_ _2779_ sg13g2_o21ai_1
Xhold307 s0.data_new_delayed\[6\] VPWR VGND net603 sg13g2_dlygate4sd3_1
X_4391_ VGND VPWR _2719_ _2716_ net1239 sg13g2_or2_1
Xhold318 _1032_ VPWR VGND net614 sg13g2_dlygate4sd3_1
X_3411_ _1835_ _1838_ net1311 _1839_ VPWR VGND sg13g2_nand3_1
X_3342_ VGND VPWR net1000 _1774_ _1775_ _1720_ sg13g2_a21oi_1
X_6130_ net145 VGND VPWR _0180_ s0.data_out\[7\]\[2\] clknet_leaf_15_clk sg13g2_dfrbpq_2
X_6061_ net219 VGND VPWR _0111_ s0.data_out\[12\]\[0\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_3273_ net991 s0.data_out\[5\]\[0\] _1714_ VPWR VGND sg13g2_and2_1
XFILLER_39_712 VPWR VGND sg13g2_fill_1
X_5012_ s0.data_out\[15\]\[0\] s0.data_out\[14\]\[0\] net1130 _0717_ VPWR VGND sg13g2_mux2_1
XFILLER_27_918 VPWR VGND sg13g2_decap_8
XFILLER_26_406 VPWR VGND sg13g2_decap_8
X_5914_ VGND VPWR net1017 net517 _1529_ _1528_ sg13g2_a21oi_1
X_5976__39 VPWR VGND net39 sg13g2_tiehi
X_5845_ VGND VPWR _2449_ net1021 _1469_ _1468_ sg13g2_a21oi_1
XFILLER_21_122 VPWR VGND sg13g2_fill_1
X_5776_ net1343 VPWR _1404_ VGND net920 _1403_ sg13g2_o21ai_1
X_4727_ VGND VPWR net1147 net456 _0459_ _0458_ sg13g2_a21oi_1
X_4658_ s0.data_out\[18\]\[4\] s0.data_out\[17\]\[4\] net1163 _0399_ VPWR VGND sg13g2_mux2_1
X_3609_ _2018_ _2017_ net1263 _2002_ net1269 VPWR VGND sg13g2_a22oi_1
X_4589_ net1158 s0.data_out\[17\]\[4\] _0334_ VPWR VGND sg13g2_and2_1
XFILLER_27_1016 VPWR VGND sg13g2_decap_8
XFILLER_27_1027 VPWR VGND sg13g2_fill_2
XFILLER_29_211 VPWR VGND sg13g2_decap_8
XFILLER_45_704 VPWR VGND sg13g2_decap_8
XFILLER_29_266 VPWR VGND sg13g2_decap_4
XFILLER_44_236 VPWR VGND sg13g2_fill_2
XFILLER_13_601 VPWR VGND sg13g2_decap_4
XFILLER_41_954 VPWR VGND sg13g2_decap_8
XFILLER_8_126 VPWR VGND sg13g2_fill_1
XFILLER_32_62 VPWR VGND sg13g2_decap_8
XFILLER_5_811 VPWR VGND sg13g2_decap_8
XFILLER_5_888 VPWR VGND sg13g2_decap_8
XFILLER_48_520 VPWR VGND sg13g2_decap_8
XFILLER_0_593 VPWR VGND sg13g2_decap_8
XFILLER_35_214 VPWR VGND sg13g2_decap_8
X_3960_ net945 net1049 _2335_ VPWR VGND sg13g2_nor2b_1
XFILLER_35_258 VPWR VGND sg13g2_fill_1
XFILLER_17_984 VPWR VGND sg13g2_decap_8
X_5966__50 VPWR VGND net50 sg13g2_tiehi
X_3891_ _2273_ _2274_ _2275_ _2276_ VPWR VGND sg13g2_nor3_1
X_5630_ net1082 VPWR _1278_ VGND _1276_ _1277_ sg13g2_o21ai_1
XFILLER_31_486 VPWR VGND sg13g2_decap_4
X_6140__134 VPWR VGND net134 sg13g2_tiehi
X_5561_ _1218_ _1217_ net1252 _1213_ net1256 VPWR VGND sg13g2_a22oi_1
X_4512_ VGND VPWR net1183 _2827_ _2828_ _2798_ sg13g2_a21oi_1
X_5492_ _1153_ net429 net1097 VPWR VGND sg13g2_nand2b_1
Xhold115 s0.data_out\[7\]\[4\] VPWR VGND net411 sg13g2_dlygate4sd3_1
Xhold126 s0.data_out\[16\]\[2\] VPWR VGND net422 sg13g2_dlygate4sd3_1
Xhold104 s0.data_out\[9\]\[3\] VPWR VGND net400 sg13g2_dlygate4sd3_1
X_4443_ net1168 net1065 _2765_ VPWR VGND sg13g2_nor2b_1
Xhold159 s0.data_out\[20\]\[1\] VPWR VGND net455 sg13g2_dlygate4sd3_1
Xhold137 s0.data_out\[4\]\[1\] VPWR VGND net433 sg13g2_dlygate4sd3_1
Xhold148 _1978_ VPWR VGND net444 sg13g2_dlygate4sd3_1
X_4374_ _2692_ VPWR _2702_ VGND net1273 _2697_ sg13g2_o21ai_1
X_6113_ net164 VGND VPWR _0163_ s0.genblk1\[8\].modules.bubble clknet_leaf_17_clk
+ sg13g2_dfrbpq_1
X_3325_ _1759_ VPWR _1760_ VGND _1755_ _1758_ sg13g2_o21ai_1
X_3256_ net313 net1209 _1701_ VPWR VGND sg13g2_nor2_1
X_6044_ net238 VGND VPWR _0094_ s0.data_out\[14\]\[7\] clknet_leaf_29_clk sg13g2_dfrbpq_2
XFILLER_39_531 VPWR VGND sg13g2_decap_8
X_3187_ _1634_ VPWR _1635_ VGND _1630_ _1633_ sg13g2_o21ai_1
XFILLER_27_726 VPWR VGND sg13g2_fill_1
XFILLER_26_214 VPWR VGND sg13g2_decap_4
XFILLER_27_737 VPWR VGND sg13g2_fill_1
XFILLER_26_247 VPWR VGND sg13g2_decap_8
X_5828_ _1394_ _1453_ net1252 _1454_ VPWR VGND sg13g2_nand3_1
X_5759_ net1027 net1059 _1389_ VPWR VGND sg13g2_nor2b_1
XFILLER_2_847 VPWR VGND sg13g2_decap_8
XFILLER_49_339 VPWR VGND sg13g2_fill_1
XFILLER_18_715 VPWR VGND sg13g2_decap_4
XFILLER_45_567 VPWR VGND sg13g2_fill_2
XFILLER_27_84 VPWR VGND sg13g2_fill_1
XFILLER_14_954 VPWR VGND sg13g2_decap_8
XFILLER_43_83 VPWR VGND sg13g2_decap_8
XFILLER_41_762 VPWR VGND sg13g2_fill_1
XFILLER_9_413 VPWR VGND sg13g2_decap_4
XFILLER_43_94 VPWR VGND sg13g2_fill_1
XFILLER_40_283 VPWR VGND sg13g2_decap_8
XFILLER_4_22 VPWR VGND sg13g2_fill_1
XFILLER_4_55 VPWR VGND sg13g2_decap_4
X_3110_ _1567_ net1025 _1566_ VPWR VGND sg13g2_nand2b_1
X_4090_ net1228 _2449_ VPWR VGND sg13g2_inv_4
XFILLER_49_884 VPWR VGND sg13g2_decap_8
X_4992_ _0698_ VPWR _0699_ VGND _0694_ _0697_ sg13g2_o21ai_1
XFILLER_23_217 VPWR VGND sg13g2_decap_8
X_3943_ _2320_ net929 _2319_ VPWR VGND sg13g2_nand2_1
XFILLER_23_239 VPWR VGND sg13g2_fill_1
X_3874_ VGND VPWR net962 _2258_ _2259_ _2219_ sg13g2_a21oi_1
XFILLER_17_1026 VPWR VGND sg13g2_fill_2
X_5613_ net1036 net1062 _1263_ VPWR VGND sg13g2_nor2b_1
Xclkbuf_3_2__f_clk clknet_0_clk clknet_3_2__leaf_clk VPWR VGND sg13g2_buf_8
X_5544_ _1200_ net1080 _1176_ _1201_ VPWR VGND sg13g2_a21o_1
X_5475_ VPWR _0124_ _1138_ VGND sg13g2_inv_1
X_4426_ net1167 s0.data_out\[18\]\[0\] _2750_ VPWR VGND sg13g2_and2_1
XFILLER_48_39 VPWR VGND sg13g2_fill_1
XFILLER_48_28 VPWR VGND sg13g2_decap_8
X_4357_ net1286 VPWR _2686_ VGND net931 _2685_ sg13g2_o21ai_1
X_4288_ _2625_ VPWR _2626_ VGND net1197 _2504_ sg13g2_o21ai_1
X_3308_ _1741_ _1744_ net1326 _1745_ VPWR VGND sg13g2_nand3_1
X_3239_ s0.data_out\[7\]\[7\] s0.data_out\[6\]\[7\] net1010 _1684_ VPWR VGND sg13g2_mux2_1
XFILLER_39_350 VPWR VGND sg13g2_decap_8
X_6027_ net256 VGND VPWR _0077_ s0.data_out\[15\]\[2\] clknet_leaf_30_clk sg13g2_dfrbpq_2
XFILLER_27_501 VPWR VGND sg13g2_decap_4
XFILLER_14_217 VPWR VGND sg13g2_decap_8
XFILLER_23_773 VPWR VGND sg13g2_fill_2
XFILLER_11_946 VPWR VGND sg13g2_decap_8
X_6201__68 VPWR VGND net68 sg13g2_tiehi
XFILLER_13_86 VPWR VGND sg13g2_fill_2
XFILLER_2_622 VPWR VGND sg13g2_decap_8
XFILLER_1_121 VPWR VGND sg13g2_decap_8
Xfanout970 net975 net970 VPWR VGND sg13g2_buf_2
XFILLER_46_810 VPWR VGND sg13g2_decap_8
XFILLER_37_309 VPWR VGND sg13g2_fill_2
Xfanout981 net982 net981 VPWR VGND sg13g2_buf_8
Xfanout992 net993 net992 VPWR VGND sg13g2_buf_8
XFILLER_46_887 VPWR VGND sg13g2_decap_8
XFILLER_33_504 VPWR VGND sg13g2_fill_2
XFILLER_33_537 VPWR VGND sg13g2_decap_8
XFILLER_41_570 VPWR VGND sg13g2_decap_8
XFILLER_9_243 VPWR VGND sg13g2_fill_2
X_3590_ VPWR _0221_ _1999_ VGND sg13g2_inv_1
X_5951__67 VPWR VGND net67 sg13g2_tiehi
Xclkload13 VPWR clkload13/Y clknet_leaf_15_clk VGND sg13g2_inv_1
XFILLER_6_961 VPWR VGND sg13g2_decap_8
X_5260_ VGND VPWR _0942_ net584 net1338 sg13g2_or2_1
X_4211_ net1204 _2552_ _2553_ _2554_ VPWR VGND sg13g2_nor3_1
X_5191_ _0880_ _0881_ _0882_ VPWR VGND sg13g2_nor2_1
X_4142_ _2498_ net1260 net912 VPWR VGND sg13g2_nand2_1
X_4073_ _2433_ VPWR _2434_ VGND net1260 _2412_ sg13g2_o21ai_1
XFILLER_49_681 VPWR VGND sg13g2_decap_8
XFILLER_37_843 VPWR VGND sg13g2_fill_1
XFILLER_37_821 VPWR VGND sg13g2_fill_1
XFILLER_37_865 VPWR VGND sg13g2_fill_1
X_4975_ _0680_ _0683_ net1322 _0684_ VPWR VGND sg13g2_nand3_1
X_3926_ s0.data_out\[0\]\[2\] s0.data_out\[1\]\[2\] net955 _2305_ VPWR VGND sg13g2_mux2_1
Xclkload7 VPWR clkload7/Y clknet_leaf_14_clk VGND sg13g2_inv_1
X_3857_ _2242_ net961 _2241_ VPWR VGND sg13g2_nand2b_1
X_3788_ _2177_ _2180_ net1297 _2181_ VPWR VGND sg13g2_nand3_1
XFILLER_30_1023 VPWR VGND sg13g2_decap_4
X_5527_ VGND VPWR net1095 _1183_ _1184_ _1140_ sg13g2_a21oi_1
X_5458_ _1123_ _1124_ _0121_ VPWR VGND sg13g2_nor2_1
XFILLER_8_1013 VPWR VGND sg13g2_decap_8
X_4409_ VPWR VGND _2720_ _2626_ _2735_ _2708_ _2737_ _2733_ sg13g2_a221oi_1
X_5389_ net1336 VPWR _1059_ VGND _2451_ _1058_ sg13g2_o21ai_1
Xfanout1209 net1210 net1209 VPWR VGND sg13g2_buf_8
XFILLER_27_342 VPWR VGND sg13g2_decap_4
XFILLER_15_559 VPWR VGND sg13g2_fill_1
XFILLER_42_356 VPWR VGND sg13g2_fill_2
XFILLER_23_581 VPWR VGND sg13g2_fill_1
XFILLER_11_754 VPWR VGND sg13g2_decap_8
XFILLER_6_246 VPWR VGND sg13g2_decap_8
XFILLER_40_95 VPWR VGND sg13g2_fill_2
XFILLER_3_964 VPWR VGND sg13g2_decap_8
Xheichips25_top_sorter_16 VPWR VGND uio_out[0] sg13g2_tielo
XFILLER_46_684 VPWR VGND sg13g2_decap_8
XFILLER_33_323 VPWR VGND sg13g2_decap_8
X_4760_ _0489_ net1152 net550 VPWR VGND sg13g2_nand2_1
X_3711_ VPWR _0232_ _2109_ VGND sg13g2_inv_1
X_4691_ VPWR _0051_ _0427_ VGND sg13g2_inv_1
X_3642_ VGND VPWR _2045_ _2049_ _0222_ _2050_ sg13g2_a21oi_1
X_3573_ _1984_ VPWR _1985_ VGND net1313 net470 sg13g2_o21ai_1
X_5312_ _0987_ VPWR _0993_ VGND _0982_ _0988_ sg13g2_o21ai_1
XFILLER_46_0 VPWR VGND sg13g2_fill_2
X_5243_ net1338 VPWR _0927_ VGND net936 _0926_ sg13g2_o21ai_1
Xhold19 s0.genblk1\[10\].modules.bubble VPWR VGND net315 sg13g2_dlygate4sd3_1
X_5174_ VGND VPWR _0867_ _0865_ net1251 sg13g2_or2_1
X_4125_ _2484_ net493 VPWR VGND sg13g2_inv_2
X_4056_ VGND VPWR net1294 _2419_ _0267_ _2417_ sg13g2_a21oi_1
XFILLER_12_518 VPWR VGND sg13g2_decap_4
X_4958_ net1138 VPWR _0669_ VGND _0667_ _0668_ sg13g2_o21ai_1
X_3909_ net1299 _2285_ _0249_ VPWR VGND sg13g2_and2_1
X_4889_ _0605_ net1135 _0558_ _0606_ VPWR VGND sg13g2_a21o_1
XFILLER_10_43 VPWR VGND sg13g2_fill_2
XFILLER_0_901 VPWR VGND sg13g2_decap_8
XFILLER_10_76 VPWR VGND sg13g2_fill_2
Xfanout1006 net1007 net1006 VPWR VGND sg13g2_buf_1
Xfanout1017 net1018 net1017 VPWR VGND sg13g2_buf_1
Xfanout1028 net1029 net1028 VPWR VGND sg13g2_buf_1
XFILLER_48_927 VPWR VGND sg13g2_decap_8
XFILLER_0_978 VPWR VGND sg13g2_decap_8
Xfanout1039 net1040 net1039 VPWR VGND sg13g2_buf_1
XFILLER_19_106 VPWR VGND sg13g2_decap_8
XFILLER_43_632 VPWR VGND sg13g2_fill_1
XFILLER_43_621 VPWR VGND sg13g2_decap_8
XFILLER_15_312 VPWR VGND sg13g2_fill_1
XFILLER_27_183 VPWR VGND sg13g2_decap_4
XFILLER_42_142 VPWR VGND sg13g2_fill_1
XFILLER_31_827 VPWR VGND sg13g2_fill_1
XFILLER_35_62 VPWR VGND sg13g2_decap_4
XFILLER_7_533 VPWR VGND sg13g2_fill_1
XFILLER_11_584 VPWR VGND sg13g2_decap_4
XFILLER_7_544 VPWR VGND sg13g2_fill_2
XFILLER_3_761 VPWR VGND sg13g2_decap_8
X_5988__26 VPWR VGND net26 sg13g2_tiehi
XFILLER_20_1011 VPWR VGND sg13g2_decap_8
XFILLER_46_470 VPWR VGND sg13g2_decap_4
X_5930_ _1536_ VPWR _1544_ VGND net1278 _1539_ sg13g2_o21ai_1
XFILLER_33_120 VPWR VGND sg13g2_decap_4
X_5861_ _1482_ VPWR _1483_ VGND net1328 net390 sg13g2_o21ai_1
XFILLER_34_687 VPWR VGND sg13g2_fill_2
X_4812_ net1134 s0.data_out\[15\]\[0\] _0537_ VPWR VGND sg13g2_and2_1
X_5792_ _1418_ net1031 net526 VPWR VGND sg13g2_nand2_1
X_4743_ VGND VPWR net1145 net591 _0473_ _0472_ sg13g2_a21oi_1
XFILLER_21_359 VPWR VGND sg13g2_fill_1
XFILLER_30_893 VPWR VGND sg13g2_fill_2
X_4674_ VGND VPWR net1222 net1151 _0413_ _0412_ sg13g2_a21oi_1
X_3625_ VGND VPWR net972 _2033_ _2034_ _1982_ sg13g2_a21oi_1
X_3556_ _1966_ _1969_ net1312 _1970_ VPWR VGND sg13g2_nand3_1
X_3487_ s0.data_out\[5\]\[6\] s0.data_out\[4\]\[6\] net988 _1908_ VPWR VGND sg13g2_mux2_1
X_5226_ VGND VPWR net1101 net472 _0912_ _0911_ sg13g2_a21oi_1
X_5157_ _0850_ net1121 net597 VPWR VGND sg13g2_nand2_1
X_4108_ VPWR _2467_ net1025 VGND sg13g2_inv_1
X_5088_ net1112 net1066 _0787_ VPWR VGND sg13g2_nor2b_1
XFILLER_38_982 VPWR VGND sg13g2_decap_8
X_4039_ net1292 net345 _2406_ VPWR VGND sg13g2_nor2_1
XFILLER_40_679 VPWR VGND sg13g2_decap_8
XFILLER_21_64 VPWR VGND sg13g2_decap_8
XFILLER_48_724 VPWR VGND sg13g2_decap_8
XFILLER_0_775 VPWR VGND sg13g2_decap_8
XFILLER_35_418 VPWR VGND sg13g2_decap_8
XFILLER_46_94 VPWR VGND sg13g2_decap_8
XFILLER_46_83 VPWR VGND sg13g2_fill_2
XFILLER_44_941 VPWR VGND sg13g2_decap_8
XFILLER_30_112 VPWR VGND sg13g2_fill_2
XFILLER_31_613 VPWR VGND sg13g2_fill_1
XFILLER_30_156 VPWR VGND sg13g2_fill_2
XFILLER_8_886 VPWR VGND sg13g2_decap_8
XFILLER_7_363 VPWR VGND sg13g2_fill_1
XFILLER_7_352 VPWR VGND sg13g2_decap_8
Xhold308 s0.data_new_delayed\[3\] VPWR VGND net604 sg13g2_dlygate4sd3_1
X_4390_ VGND VPWR _2718_ _2712_ net1231 sg13g2_or2_1
X_3410_ net990 VPWR _1838_ VGND _1836_ _1837_ sg13g2_o21ai_1
X_3341_ _1773_ net991 _1721_ _1774_ VPWR VGND sg13g2_a21o_1
X_6060_ net220 VGND VPWR _0110_ s0.valid_out\[12\][0] clknet_leaf_27_clk sg13g2_dfrbpq_2
X_3272_ _1713_ net916 _1712_ VPWR VGND sg13g2_nand2_1
X_5011_ _0659_ _0715_ _0716_ VPWR VGND sg13g2_and2_1
XFILLER_39_746 VPWR VGND sg13g2_decap_8
XFILLER_38_278 VPWR VGND sg13g2_decap_8
X_5913_ net1017 net1048 _1528_ VPWR VGND sg13g2_nor2b_1
XFILLER_35_985 VPWR VGND sg13g2_decap_8
X_5844_ net1025 VPWR _1468_ VGND net1230 net1016 sg13g2_o21ai_1
XFILLER_22_657 VPWR VGND sg13g2_fill_1
X_5775_ VGND VPWR net1027 s0.data_out\[8\]\[6\] _1403_ _1402_ sg13g2_a21oi_1
X_4726_ net1146 net1053 _0458_ VPWR VGND sg13g2_nor2b_1
X_4657_ _0397_ VPWR _0398_ VGND net1262 _0378_ sg13g2_o21ai_1
X_3608_ _1966_ _2016_ _2017_ VPWR VGND sg13g2_and2_1
X_4588_ _0333_ net925 _0332_ VPWR VGND sg13g2_nand2_1
X_3539_ net980 VPWR _1955_ VGND _1953_ _1954_ sg13g2_o21ai_1
X_5209_ net1100 s0.data_out\[12\]\[1\] _0897_ VPWR VGND sg13g2_and2_1
X_6189_ net81 VGND VPWR _0239_ s0.data_out\[2\]\[1\] clknet_leaf_6_clk sg13g2_dfrbpq_2
XFILLER_29_245 VPWR VGND sg13g2_fill_1
XFILLER_44_204 VPWR VGND sg13g2_fill_2
XFILLER_26_930 VPWR VGND sg13g2_fill_1
XFILLER_16_53 VPWR VGND sg13g2_decap_4
XFILLER_41_933 VPWR VGND sg13g2_decap_8
XFILLER_16_75 VPWR VGND sg13g2_fill_1
XFILLER_8_138 VPWR VGND sg13g2_fill_1
XFILLER_10_1010 VPWR VGND sg13g2_decap_8
XFILLER_5_867 VPWR VGND sg13g2_decap_8
XFILLER_4_377 VPWR VGND sg13g2_fill_1
X_6133__142 VPWR VGND net142 sg13g2_tiehi
XFILLER_0_572 VPWR VGND sg13g2_decap_8
XFILLER_36_716 VPWR VGND sg13g2_decap_8
XFILLER_48_598 VPWR VGND sg13g2_decap_8
XFILLER_17_963 VPWR VGND sg13g2_decap_8
XFILLER_43_292 VPWR VGND sg13g2_decap_4
XFILLER_43_281 VPWR VGND sg13g2_fill_2
X_3890_ _2275_ net1214 _2267_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_421 VPWR VGND sg13g2_decap_4
XFILLER_31_454 VPWR VGND sg13g2_decap_4
X_5560_ VGND VPWR net1093 _1216_ _1217_ _1161_ sg13g2_a21oi_1
X_4511_ _2826_ net1168 _2799_ _2827_ VPWR VGND sg13g2_a21o_1
X_5491_ VPWR _0126_ _1152_ VGND sg13g2_inv_1
XFILLER_7_171 VPWR VGND sg13g2_fill_1
X_4442_ net1167 s0.data_out\[18\]\[2\] _2764_ VPWR VGND sg13g2_and2_1
Xhold105 s0.data_out\[17\]\[4\] VPWR VGND net401 sg13g2_dlygate4sd3_1
Xhold116 s0.data_out\[6\]\[0\] VPWR VGND net412 sg13g2_dlygate4sd3_1
Xhold138 s0.data_out\[8\]\[3\] VPWR VGND net434 sg13g2_dlygate4sd3_1
Xhold149 s0.data_out\[15\]\[2\] VPWR VGND net445 sg13g2_dlygate4sd3_1
Xhold127 s0.data_out\[6\]\[4\] VPWR VGND net423 sg13g2_dlygate4sd3_1
X_4373_ VPWR VGND _2634_ net1281 _2700_ net1273 _2701_ _2697_ sg13g2_a221oi_1
X_3324_ VGND VPWR _1759_ net557 net1325 sg13g2_or2_1
X_6112_ net165 VGND VPWR _0162_ s0.shift_out\[9\][0] clknet_leaf_19_clk sg13g2_dfrbpq_2
XFILLER_39_510 VPWR VGND sg13g2_decap_8
X_3255_ _1699_ VPWR _1700_ VGND _1682_ _1696_ sg13g2_o21ai_1
X_6043_ net239 VGND VPWR _0093_ s0.data_out\[14\]\[6\] clknet_leaf_31_clk sg13g2_dfrbpq_2
X_3186_ VGND VPWR _1634_ net589 net1329 sg13g2_or2_1
XFILLER_2_1008 VPWR VGND sg13g2_decap_8
XFILLER_26_204 VPWR VGND sg13g2_fill_1
X_5827_ _1453_ net1037 _1452_ VPWR VGND sg13g2_nand2b_1
XFILLER_23_999 VPWR VGND sg13g2_decap_8
X_5758_ net1027 s0.data_out\[8\]\[4\] _1388_ VPWR VGND sg13g2_and2_1
X_4709_ _0443_ net924 _0442_ VPWR VGND sg13g2_nand2_1
X_5689_ _1334_ net1082 _1333_ VPWR VGND sg13g2_nand2b_1
XFILLER_2_826 VPWR VGND sg13g2_decap_8
XFILLER_49_318 VPWR VGND sg13g2_decap_8
X_6117__159 VPWR VGND net159 sg13g2_tiehi
XFILLER_17_204 VPWR VGND sg13g2_fill_2
XFILLER_27_41 VPWR VGND sg13g2_fill_1
XFILLER_27_52 VPWR VGND sg13g2_decap_8
XFILLER_45_557 VPWR VGND sg13g2_fill_1
XFILLER_27_96 VPWR VGND sg13g2_fill_1
XFILLER_33_719 VPWR VGND sg13g2_decap_4
XFILLER_32_229 VPWR VGND sg13g2_decap_8
XFILLER_9_403 VPWR VGND sg13g2_fill_2
X_5963__54 VPWR VGND net54 sg13g2_tiehi
XFILLER_4_141 VPWR VGND sg13g2_decap_4
XFILLER_4_152 VPWR VGND sg13g2_decap_8
XFILLER_4_78 VPWR VGND sg13g2_decap_8
XFILLER_49_863 VPWR VGND sg13g2_decap_8
X_4991_ VGND VPWR _0698_ net562 net1319 sg13g2_or2_1
X_3942_ s0.data_out\[0\]\[4\] s0.data_out\[1\]\[4\] net956 _2319_ VPWR VGND sg13g2_mux2_1
XFILLER_17_1005 VPWR VGND sg13g2_decap_8
XFILLER_32_741 VPWR VGND sg13g2_fill_1
X_3873_ _2257_ net954 _2220_ _2258_ VPWR VGND sg13g2_a21o_1
XFILLER_20_914 VPWR VGND sg13g2_fill_1
XFILLER_31_284 VPWR VGND sg13g2_fill_1
X_5612_ net1036 s0.data_out\[9\]\[3\] _1262_ VPWR VGND sg13g2_and2_1
X_5543_ s0.data_out\[11\]\[7\] s0.data_out\[10\]\[7\] net1085 _1200_ VPWR VGND sg13g2_mux2_1
XFILLER_9_992 VPWR VGND sg13g2_decap_8
X_5474_ _1137_ VPWR _1138_ VGND _1133_ _1136_ sg13g2_o21ai_1
X_4425_ _2749_ net926 _2748_ VPWR VGND sg13g2_nand2_1
X_4356_ VGND VPWR net1180 s0.data_out\[19\]\[7\] _2685_ _2684_ sg13g2_a21oi_1
X_3307_ net1000 VPWR _1744_ VGND _1742_ _1743_ sg13g2_o21ai_1
X_4287_ _2625_ _2624_ _2623_ VPWR VGND sg13g2_nand2b_1
X_3238_ _1683_ net1009 net519 VPWR VGND sg13g2_nand2_1
X_6026_ net257 VGND VPWR _0076_ s0.data_out\[15\]\[1\] clknet_leaf_30_clk sg13g2_dfrbpq_2
X_3169_ net1327 VPWR _1619_ VGND net917 _1618_ sg13g2_o21ai_1
XFILLER_27_557 VPWR VGND sg13g2_decap_4
XFILLER_27_568 VPWR VGND sg13g2_fill_2
XFILLER_14_207 VPWR VGND sg13g2_fill_1
XFILLER_22_273 VPWR VGND sg13g2_decap_8
XFILLER_7_929 VPWR VGND sg13g2_decap_8
X_5960__57 VPWR VGND net57 sg13g2_tiehi
XFILLER_2_601 VPWR VGND sg13g2_decap_8
XFILLER_1_166 VPWR VGND sg13g2_fill_2
XFILLER_49_126 VPWR VGND sg13g2_decap_4
Xfanout960 s0.shift_out\[2\][0] net960 VPWR VGND sg13g2_buf_8
XFILLER_38_40 VPWR VGND sg13g2_fill_2
Xfanout971 net975 net971 VPWR VGND sg13g2_buf_8
Xfanout993 s0.shift_out\[5\][0] net993 VPWR VGND sg13g2_buf_2
Xfanout982 net986 net982 VPWR VGND sg13g2_buf_8
X_6130__145 VPWR VGND net145 sg13g2_tiehi
XFILLER_46_866 VPWR VGND sg13g2_decap_8
XFILLER_18_546 VPWR VGND sg13g2_fill_1
XFILLER_14_741 VPWR VGND sg13g2_decap_8
XFILLER_26_590 VPWR VGND sg13g2_decap_4
XFILLER_14_752 VPWR VGND sg13g2_fill_1
Xclkload14 VPWR clkload14/Y clknet_leaf_16_clk VGND sg13g2_inv_1
XFILLER_6_940 VPWR VGND sg13g2_decap_8
X_4210_ s0.valid_out\[21\][0] s0.data_out\[20\]\[5\] _2553_ VPWR VGND sg13g2_nor2_1
X_5190_ VGND VPWR _2449_ net1119 _0881_ net1114 sg13g2_a21oi_1
X_4141_ VGND VPWR net1211 net913 net4 _2497_ sg13g2_a21oi_1
XFILLER_49_660 VPWR VGND sg13g2_decap_8
XFILLER_23_1020 VPWR VGND sg13g2_decap_8
X_4072_ _2433_ net1214 _2414_ VPWR VGND sg13g2_nand2b_1
XFILLER_36_310 VPWR VGND sg13g2_decap_8
XFILLER_36_321 VPWR VGND sg13g2_fill_2
XFILLER_24_527 VPWR VGND sg13g2_decap_8
X_4974_ net1139 VPWR _0683_ VGND _0681_ _0682_ sg13g2_o21ai_1
X_3925_ VPWR _0251_ net397 VGND sg13g2_inv_1
Xclkload8 VPWR clkload8/Y clknet_leaf_30_clk VGND sg13g2_inv_1
X_3856_ VGND VPWR net950 _2240_ _2241_ _2179_ sg13g2_a21oi_1
X_3787_ net961 VPWR _2180_ VGND _2178_ _2179_ sg13g2_o21ai_1
XFILLER_30_1002 VPWR VGND sg13g2_decap_8
X_6077__202 VPWR VGND net202 sg13g2_tiehi
X_5526_ _1182_ net1078 _1141_ _1183_ VPWR VGND sg13g2_a21o_1
X_5457_ net1336 VPWR _1124_ VGND net413 _1119_ sg13g2_o21ai_1
X_4408_ _2736_ _2718_ _2717_ VPWR VGND sg13g2_nand2b_1
X_5388_ VGND VPWR net1091 net540 _1058_ _1057_ sg13g2_a21oi_1
X_4339_ net1183 s0.data_out\[19\]\[5\] _2670_ VPWR VGND sg13g2_and2_1
XFILLER_47_619 VPWR VGND sg13g2_decap_8
X_6009_ net276 VGND VPWR _0059_ s0.shift_out\[17\][0] clknet_leaf_33_clk sg13g2_dfrbpq_1
XFILLER_28_844 VPWR VGND sg13g2_fill_1
XFILLER_43_825 VPWR VGND sg13g2_decap_4
XFILLER_11_733 VPWR VGND sg13g2_decap_8
XFILLER_6_214 VPWR VGND sg13g2_decap_8
XFILLER_40_30 VPWR VGND sg13g2_fill_1
XFILLER_3_943 VPWR VGND sg13g2_decap_8
XFILLER_2_431 VPWR VGND sg13g2_decap_8
XFILLER_46_1020 VPWR VGND sg13g2_decap_8
XFILLER_2_464 VPWR VGND sg13g2_decap_4
XFILLER_49_61 VPWR VGND sg13g2_fill_1
XFILLER_37_118 VPWR VGND sg13g2_decap_4
XFILLER_1_35 VPWR VGND sg13g2_decap_4
XFILLER_46_641 VPWR VGND sg13g2_decap_8
Xheichips25_top_sorter_17 VPWR VGND uio_out[1] sg13g2_tielo
XFILLER_19_844 VPWR VGND sg13g2_fill_2
XFILLER_46_663 VPWR VGND sg13g2_decap_8
XFILLER_33_302 VPWR VGND sg13g2_fill_2
X_3710_ _2108_ VPWR _2109_ VGND _2104_ _2107_ sg13g2_o21ai_1
XFILLER_42_880 VPWR VGND sg13g2_decap_8
X_4690_ _0426_ VPWR _0427_ VGND net1304 net468 sg13g2_o21ai_1
X_3641_ VGND VPWR _2050_ net1210 net317 sg13g2_or2_1
X_3572_ _1980_ _1983_ net1313 _1984_ VPWR VGND sg13g2_nand3_1
X_5311_ _0992_ _0977_ _0987_ _0991_ VPWR VGND sg13g2_and3_1
X_5242_ VGND VPWR net1106 net501 _0926_ _0925_ sg13g2_a21oi_1
XFILLER_39_0 VPWR VGND sg13g2_fill_2
X_5173_ net1251 _0865_ _0866_ VPWR VGND sg13g2_nor2_1
X_4124_ VPWR _2483_ s0.data_out\[19\]\[2\] VGND sg13g2_inv_1
X_4055_ _2418_ VPWR _2419_ VGND _2465_ net1053 sg13g2_o21ai_1
XFILLER_24_335 VPWR VGND sg13g2_fill_1
X_4957_ net1122 net1066 _0668_ VPWR VGND sg13g2_nor2b_1
X_3908_ VGND VPWR _2442_ _2285_ _0248_ _2290_ sg13g2_a21oi_1
X_4888_ _0604_ VPWR _0605_ VGND net1141 _2485_ sg13g2_o21ai_1
X_3839_ _2225_ net495 net966 VPWR VGND sg13g2_nand2b_1
XFILLER_20_596 VPWR VGND sg13g2_fill_2
X_5509_ VGND VPWR _1087_ _1167_ _1168_ net1093 sg13g2_a21oi_1
Xfanout1018 net339 net1018 VPWR VGND sg13g2_buf_8
Xfanout1007 s0.shift_out\[6\][0] net1007 VPWR VGND sg13g2_buf_2
Xfanout1029 s0.shift_out\[8\][0] net1029 VPWR VGND sg13g2_buf_1
XFILLER_0_957 VPWR VGND sg13g2_decap_8
XFILLER_48_906 VPWR VGND sg13g2_decap_8
XFILLER_47_449 VPWR VGND sg13g2_decap_8
XFILLER_19_75 VPWR VGND sg13g2_fill_1
XFILLER_19_86 VPWR VGND sg13g2_fill_2
XFILLER_28_652 VPWR VGND sg13g2_fill_2
XFILLER_28_674 VPWR VGND sg13g2_fill_2
XFILLER_15_335 VPWR VGND sg13g2_decap_8
XFILLER_27_195 VPWR VGND sg13g2_fill_2
XFILLER_43_677 VPWR VGND sg13g2_fill_2
XFILLER_43_688 VPWR VGND sg13g2_decap_8
XFILLER_24_891 VPWR VGND sg13g2_fill_2
XFILLER_35_96 VPWR VGND sg13g2_decap_8
XFILLER_42_198 VPWR VGND sg13g2_fill_2
XFILLER_3_740 VPWR VGND sg13g2_decap_8
XFILLER_32_7 VPWR VGND sg13g2_decap_4
XFILLER_39_906 VPWR VGND sg13g2_decap_4
XFILLER_38_405 VPWR VGND sg13g2_fill_1
XFILLER_47_983 VPWR VGND sg13g2_decap_8
X_5860_ _1478_ _1481_ net1328 _1482_ VPWR VGND sg13g2_nand3_1
X_4811_ _0536_ net922 _0535_ VPWR VGND sg13g2_nand2_1
XFILLER_21_316 VPWR VGND sg13g2_fill_1
X_5791_ _1373_ VPWR _1417_ VGND net919 _1416_ sg13g2_o21ai_1
X_4742_ net1145 net1045 _0472_ VPWR VGND sg13g2_nor2b_1
X_4673_ net1161 VPWR _0412_ VGND net1226 net1146 sg13g2_o21ai_1
X_3624_ s0.data_out\[4\]\[5\] s0.data_out\[3\]\[5\] net978 _2033_ VPWR VGND sg13g2_mux2_1
X_3555_ net980 VPWR _1969_ VGND _1967_ _1968_ sg13g2_o21ai_1
X_3486_ _1907_ net988 net511 VPWR VGND sg13g2_nand2_1
X_6074__205 VPWR VGND net205 sg13g2_tiehi
X_5225_ net1101 net1063 _0911_ VPWR VGND sg13g2_nor2b_1
XFILLER_5_1028 VPWR VGND sg13g2_fill_1
X_5156_ VGND VPWR net1128 _0848_ _0849_ _0821_ sg13g2_a21oi_1
X_5950__221 VPWR VGND net221 sg13g2_tiehi
X_4107_ VPWR _2466_ net1037 VGND sg13g2_inv_1
X_5087_ VGND VPWR _0707_ _0785_ _0786_ net1127 sg13g2_a21oi_1
XFILLER_29_449 VPWR VGND sg13g2_fill_2
XFILLER_38_961 VPWR VGND sg13g2_decap_8
X_4038_ VPWR _0263_ _2405_ VGND sg13g2_inv_1
XFILLER_37_493 VPWR VGND sg13g2_decap_8
XFILLER_24_143 VPWR VGND sg13g2_decap_4
XFILLER_40_625 VPWR VGND sg13g2_decap_4
X_5989_ net25 VGND VPWR _0039_ s0.data_out\[18\]\[0\] clknet_leaf_35_clk sg13g2_dfrbpq_2
XFILLER_12_305 VPWR VGND sg13g2_fill_1
XFILLER_24_176 VPWR VGND sg13g2_fill_2
XFILLER_25_699 VPWR VGND sg13g2_fill_2
XFILLER_12_338 VPWR VGND sg13g2_decap_8
XFILLER_21_850 VPWR VGND sg13g2_fill_2
XFILLER_21_894 VPWR VGND sg13g2_fill_2
XFILLER_21_87 VPWR VGND sg13g2_fill_1
XFILLER_21_98 VPWR VGND sg13g2_decap_8
XFILLER_48_703 VPWR VGND sg13g2_decap_8
XFILLER_0_754 VPWR VGND sg13g2_decap_8
XFILLER_46_51 VPWR VGND sg13g2_decap_8
XFILLER_44_920 VPWR VGND sg13g2_decap_8
XFILLER_16_611 VPWR VGND sg13g2_decap_4
XFILLER_44_997 VPWR VGND sg13g2_decap_8
XFILLER_43_485 VPWR VGND sg13g2_decap_8
XFILLER_15_198 VPWR VGND sg13g2_fill_1
XFILLER_7_331 VPWR VGND sg13g2_fill_1
XFILLER_7_320 VPWR VGND sg13g2_decap_8
XFILLER_12_894 VPWR VGND sg13g2_fill_1
XFILLER_7_89 VPWR VGND sg13g2_decap_8
Xhold309 s0.data_new_delayed\[1\] VPWR VGND net605 sg13g2_dlygate4sd3_1
X_3340_ s0.data_out\[6\]\[1\] s0.data_out\[5\]\[1\] net997 _1773_ VPWR VGND sg13g2_mux2_1
X_5010_ _0715_ net1138 _0714_ VPWR VGND sg13g2_nand2b_1
X_3271_ s0.data_out\[5\]\[0\] s0.data_out\[6\]\[0\] net1008 _1712_ VPWR VGND sg13g2_mux2_1
XFILLER_38_202 VPWR VGND sg13g2_decap_4
XFILLER_38_246 VPWR VGND sg13g2_fill_1
XFILLER_47_780 VPWR VGND sg13g2_decap_8
XFILLER_19_493 VPWR VGND sg13g2_decap_4
X_5912_ VGND VPWR _1436_ _1526_ _1527_ net1026 sg13g2_a21oi_1
XFILLER_35_964 VPWR VGND sg13g2_decap_8
XFILLER_34_452 VPWR VGND sg13g2_decap_4
X_5843_ net1329 net307 _0163_ VPWR VGND sg13g2_and2_1
XFILLER_22_636 VPWR VGND sg13g2_fill_2
X_5774_ net1027 net1052 _1402_ VPWR VGND sg13g2_nor2b_1
XFILLER_21_146 VPWR VGND sg13g2_fill_2
X_4725_ VGND VPWR _0393_ _0456_ _0457_ net1162 sg13g2_a21oi_1
X_4656_ _0397_ net1248 _0396_ VPWR VGND sg13g2_nand2_1
X_4587_ s0.data_out\[17\]\[4\] s0.data_out\[18\]\[4\] net1176 _0332_ VPWR VGND sg13g2_mux2_1
X_3607_ _2016_ net980 _2015_ VPWR VGND sg13g2_nand2b_1
X_3538_ net969 net1072 _1954_ VPWR VGND sg13g2_nor2b_1
XFILLER_1_529 VPWR VGND sg13g2_decap_8
X_3469_ _1890_ net990 _1889_ VPWR VGND sg13g2_nand2b_1
X_5208_ _0896_ net935 _0895_ VPWR VGND sg13g2_nand2_1
X_6188_ net82 VGND VPWR _0238_ s0.data_out\[2\]\[0\] clknet_leaf_6_clk sg13g2_dfrbpq_2
X_5139_ _0831_ net1112 _0780_ _0832_ VPWR VGND sg13g2_a21o_1
XFILLER_45_739 VPWR VGND sg13g2_decap_8
XFILLER_44_238 VPWR VGND sg13g2_fill_1
XFILLER_44_227 VPWR VGND sg13g2_fill_2
XFILLER_16_10 VPWR VGND sg13g2_decap_8
XFILLER_44_249 VPWR VGND sg13g2_decap_8
XFILLER_41_912 VPWR VGND sg13g2_decap_8
XFILLER_40_400 VPWR VGND sg13g2_decap_8
X_5975__41 VPWR VGND net41 sg13g2_tiehi
X_6126__150 VPWR VGND net150 sg13g2_tiehi
XFILLER_40_444 VPWR VGND sg13g2_fill_2
XFILLER_41_989 VPWR VGND sg13g2_decap_8
XFILLER_12_146 VPWR VGND sg13g2_fill_2
XFILLER_32_86 VPWR VGND sg13g2_decap_8
XFILLER_32_97 VPWR VGND sg13g2_fill_1
XFILLER_5_846 VPWR VGND sg13g2_decap_8
XFILLER_0_551 VPWR VGND sg13g2_decap_8
XFILLER_48_577 VPWR VGND sg13g2_decap_8
XFILLER_44_794 VPWR VGND sg13g2_decap_8
X_6209__247 VPWR VGND net247 sg13g2_tiehi
XFILLER_32_989 VPWR VGND sg13g2_decap_8
XFILLER_12_691 VPWR VGND sg13g2_fill_1
X_4510_ s0.data_out\[19\]\[7\] s0.data_out\[18\]\[7\] net1174 _2826_ VPWR VGND sg13g2_mux2_1
X_5490_ _1151_ VPWR _1152_ VGND _1147_ _1150_ sg13g2_o21ai_1
XFILLER_8_684 VPWR VGND sg13g2_fill_2
X_4441_ _2763_ net926 _2762_ VPWR VGND sg13g2_nand2_1
Xhold117 s0.was_valid_out\[11\][0] VPWR VGND net413 sg13g2_dlygate4sd3_1
Xhold106 s0.data_out\[5\]\[4\] VPWR VGND net402 sg13g2_dlygate4sd3_1
Xhold139 s0.was_valid_out\[20\][0] VPWR VGND net435 sg13g2_dlygate4sd3_1
Xhold128 s0.data_out\[2\]\[0\] VPWR VGND net424 sg13g2_dlygate4sd3_1
X_6111_ net166 VGND VPWR _0161_ s0.data_out\[9\]\[7\] clknet_leaf_19_clk sg13g2_dfrbpq_2
X_4372_ _2700_ net1193 _2699_ VPWR VGND sg13g2_nand2b_1
X_3323_ net1325 VPWR _1758_ VGND net916 _1757_ sg13g2_o21ai_1
X_3254_ VGND VPWR _1695_ _1697_ _1699_ _1698_ sg13g2_a21oi_1
X_6042_ net240 VGND VPWR _0092_ s0.data_out\[14\]\[5\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_3185_ net1326 VPWR _1633_ VGND _2468_ _1632_ sg13g2_o21ai_1
Xfanout1190 net1191 net1190 VPWR VGND sg13g2_buf_8
XFILLER_27_717 VPWR VGND sg13g2_decap_8
XFILLER_35_794 VPWR VGND sg13g2_fill_2
XFILLER_22_411 VPWR VGND sg13g2_decap_8
XFILLER_22_422 VPWR VGND sg13g2_fill_2
X_5826_ VGND VPWR net1027 _1451_ _1452_ _1396_ sg13g2_a21oi_1
XFILLER_23_978 VPWR VGND sg13g2_decap_8
XFILLER_33_1011 VPWR VGND sg13g2_decap_8
X_5757_ _1387_ net919 _1386_ VPWR VGND sg13g2_nand2_1
X_5972__44 VPWR VGND net44 sg13g2_tiehi
X_4708_ _0374_ VPWR _0442_ VGND net1164 _2485_ sg13g2_o21ai_1
X_5688_ VGND VPWR net1038 _1332_ _1333_ _1277_ sg13g2_a21oi_1
X_4639_ _0379_ VPWR _0380_ VGND _0372_ _0373_ sg13g2_o21ai_1
XFILLER_2_805 VPWR VGND sg13g2_decap_8
XFILLER_40_1015 VPWR VGND sg13g2_decap_8
XFILLER_17_216 VPWR VGND sg13g2_fill_2
XFILLER_17_238 VPWR VGND sg13g2_fill_2
XFILLER_14_901 VPWR VGND sg13g2_decap_8
XFILLER_14_912 VPWR VGND sg13g2_fill_2
XFILLER_14_923 VPWR VGND sg13g2_fill_2
XFILLER_41_786 VPWR VGND sg13g2_fill_2
XFILLER_14_989 VPWR VGND sg13g2_decap_8
XFILLER_9_459 VPWR VGND sg13g2_decap_8
XFILLER_5_610 VPWR VGND sg13g2_fill_1
XFILLER_5_687 VPWR VGND sg13g2_fill_1
XFILLER_4_13 VPWR VGND sg13g2_decap_8
XFILLER_49_842 VPWR VGND sg13g2_decap_8
XFILLER_1_893 VPWR VGND sg13g2_decap_8
XFILLER_48_363 VPWR VGND sg13g2_fill_2
XFILLER_36_525 VPWR VGND sg13g2_decap_8
XFILLER_36_569 VPWR VGND sg13g2_fill_2
X_4990_ net1320 VPWR _0697_ VGND net921 _0696_ sg13g2_o21ai_1
XFILLER_16_260 VPWR VGND sg13g2_fill_1
XFILLER_16_293 VPWR VGND sg13g2_fill_1
X_3941_ VPWR _0253_ net514 VGND sg13g2_inv_1
X_3872_ s0.data_out\[2\]\[6\] s0.data_out\[1\]\[6\] net957 _2257_ VPWR VGND sg13g2_mux2_1
XFILLER_17_1028 VPWR VGND sg13g2_fill_1
XFILLER_20_959 VPWR VGND sg13g2_decap_8
X_5611_ _1261_ net934 _1260_ VPWR VGND sg13g2_nand2_1
XFILLER_9_971 VPWR VGND sg13g2_decap_8
X_5542_ _1199_ net1085 net531 VPWR VGND sg13g2_nand2_1
X_5473_ VGND VPWR _1137_ net536 net1334 sg13g2_or2_1
X_4424_ s0.data_out\[18\]\[0\] s0.data_out\[19\]\[0\] net1187 _2748_ VPWR VGND sg13g2_mux2_1
X_4355_ net1180 net1045 _2684_ VPWR VGND sg13g2_nor2b_1
X_3306_ net992 net1059 _1743_ VPWR VGND sg13g2_nor2b_1
X_4286_ _2624_ net1222 net1189 VPWR VGND sg13g2_nand2_1
X_6116__160 VPWR VGND net160 sg13g2_tiehi
X_3237_ _1682_ _1677_ _1681_ VPWR VGND sg13g2_nand2_1
X_6025_ net258 VGND VPWR _0075_ s0.data_out\[15\]\[0\] clknet_leaf_30_clk sg13g2_dfrbpq_2
XFILLER_27_536 VPWR VGND sg13g2_decap_8
X_3168_ VGND VPWR net1002 net454 _1618_ _1617_ sg13g2_a21oi_1
XFILLER_27_547 VPWR VGND sg13g2_fill_1
XFILLER_22_252 VPWR VGND sg13g2_fill_2
XFILLER_7_908 VPWR VGND sg13g2_decap_8
X_5809_ _1433_ _1434_ _1435_ VPWR VGND _1428_ sg13g2_nand3b_1
X_6123__153 VPWR VGND net153 sg13g2_tiehi
XFILLER_13_44 VPWR VGND sg13g2_fill_1
XFILLER_13_88 VPWR VGND sg13g2_fill_1
XFILLER_8_4 VPWR VGND sg13g2_fill_1
XFILLER_49_105 VPWR VGND sg13g2_decap_8
XFILLER_2_668 VPWR VGND sg13g2_decap_8
Xfanout950 net951 net950 VPWR VGND sg13g2_buf_8
Xfanout961 s0.shift_out\[2\][0] net961 VPWR VGND sg13g2_buf_8
Xfanout994 net996 net994 VPWR VGND sg13g2_buf_8
Xfanout983 net985 net983 VPWR VGND sg13g2_buf_8
Xfanout972 net974 net972 VPWR VGND sg13g2_buf_8
XFILLER_45_311 VPWR VGND sg13g2_fill_2
XFILLER_46_845 VPWR VGND sg13g2_decap_8
XFILLER_45_366 VPWR VGND sg13g2_decap_8
XFILLER_14_797 VPWR VGND sg13g2_fill_2
Xclkload15 clknet_leaf_22_clk clkload15/Y VPWR VGND sg13g2_inv_4
XFILLER_6_996 VPWR VGND sg13g2_decap_8
XFILLER_5_462 VPWR VGND sg13g2_decap_4
X_4140_ s0.data_out\[21\]\[2\] net913 _2497_ VPWR VGND sg13g2_nor2_1
XFILLER_1_690 VPWR VGND sg13g2_decap_8
X_4071_ VPWR VGND net1260 _2431_ _2412_ net1268 _2432_ _2409_ sg13g2_a221oi_1
XFILLER_37_856 VPWR VGND sg13g2_decap_8
X_4973_ net1126 net1059 _0682_ VPWR VGND sg13g2_nor2b_1
X_3924_ _2303_ VPWR _2304_ VGND net1293 net396 sg13g2_o21ai_1
XFILLER_20_723 VPWR VGND sg13g2_decap_4
XFILLER_32_583 VPWR VGND sg13g2_decap_8
Xclkload9 clknet_leaf_31_clk clkload9/X VPWR VGND sg13g2_buf_8
X_3855_ s0.data_out\[2\]\[0\] s0.data_out\[1\]\[0\] net955 _2240_ VPWR VGND sg13g2_mux2_1
XFILLER_20_778 VPWR VGND sg13g2_fill_1
X_3786_ net949 net1073 _2179_ VPWR VGND sg13g2_nor2b_1
X_5525_ s0.data_out\[11\]\[2\] s0.data_out\[10\]\[2\] net1084 _1182_ VPWR VGND sg13g2_mux2_1
X_5456_ VGND VPWR _1117_ _1120_ _1123_ _1122_ sg13g2_a21oi_1
X_4407_ _2735_ _2728_ _2734_ VPWR VGND sg13g2_nand2_1
X_5387_ net1091 net1047 _1057_ VPWR VGND sg13g2_nor2b_1
X_4338_ _2669_ net931 _2668_ VPWR VGND sg13g2_nand2_1
X_4269_ VGND VPWR net1205 _2608_ _2609_ _2554_ sg13g2_a21oi_1
X_6008_ net277 VGND VPWR _0058_ s0.data_out\[17\]\[7\] clknet_leaf_33_clk sg13g2_dfrbpq_2
XFILLER_27_322 VPWR VGND sg13g2_fill_1
XFILLER_27_333 VPWR VGND sg13g2_decap_4
XFILLER_27_377 VPWR VGND sg13g2_fill_1
XFILLER_28_889 VPWR VGND sg13g2_decap_4
XFILLER_24_10 VPWR VGND sg13g2_decap_8
XFILLER_24_21 VPWR VGND sg13g2_fill_2
XFILLER_24_87 VPWR VGND sg13g2_fill_1
XFILLER_3_922 VPWR VGND sg13g2_decap_8
XFILLER_3_999 VPWR VGND sg13g2_decap_8
XFILLER_49_51 VPWR VGND sg13g2_fill_1
XFILLER_18_300 VPWR VGND sg13g2_decap_8
XFILLER_19_812 VPWR VGND sg13g2_fill_2
XFILLER_19_823 VPWR VGND sg13g2_decap_4
XFILLER_46_631 VPWR VGND sg13g2_fill_1
XFILLER_46_620 VPWR VGND sg13g2_decap_8
Xheichips25_top_sorter_18 VPWR VGND uio_out[3] sg13g2_tielo
XFILLER_18_311 VPWR VGND sg13g2_fill_1
XFILLER_34_837 VPWR VGND sg13g2_decap_8
XFILLER_14_572 VPWR VGND sg13g2_fill_2
XFILLER_41_391 VPWR VGND sg13g2_decap_4
X_3640_ _2047_ _2048_ _2049_ VPWR VGND sg13g2_and2_1
X_3571_ net983 VPWR _1983_ VGND _1981_ _1982_ sg13g2_o21ai_1
X_5310_ _0988_ _0989_ _0990_ _0991_ VPWR VGND sg13g2_nor3_1
XFILLER_46_2 VPWR VGND sg13g2_fill_1
X_5241_ net1106 net1056 _0925_ VPWR VGND sg13g2_nor2b_1
X_5172_ VGND VPWR net1129 _0864_ _0865_ _0807_ sg13g2_a21oi_1
X_4123_ VPWR _2482_ net368 VGND sg13g2_inv_1
X_4054_ net344 net947 net944 _2418_ VPWR VGND sg13g2_a21o_1
XFILLER_37_631 VPWR VGND sg13g2_decap_4
XFILLER_37_664 VPWR VGND sg13g2_fill_2
XFILLER_37_697 VPWR VGND sg13g2_decap_4
X_4956_ net1122 s0.data_out\[14\]\[2\] _0667_ VPWR VGND sg13g2_and2_1
X_3907_ net1298 VPWR _2290_ VGND _2287_ _2289_ sg13g2_o21ai_1
X_4887_ _0604_ net1141 net387 VPWR VGND sg13g2_nand2_1
X_3838_ VPWR _0244_ net492 VGND sg13g2_inv_1
X_6120__156 VPWR VGND net156 sg13g2_tiehi
X_3769_ VGND VPWR _2161_ _2164_ _0234_ _2165_ sg13g2_a21oi_1
XFILLER_4_719 VPWR VGND sg13g2_decap_4
X_5508_ _1167_ net521 net1097 VPWR VGND sg13g2_nand2b_1
X_5439_ _1105_ _1106_ _1104_ _1108_ VPWR VGND sg13g2_nand3_1
Xfanout1019 net1022 net1019 VPWR VGND sg13g2_buf_8
XFILLER_0_936 VPWR VGND sg13g2_decap_8
Xfanout1008 net1011 net1008 VPWR VGND sg13g2_buf_8
XFILLER_19_43 VPWR VGND sg13g2_decap_8
XFILLER_15_303 VPWR VGND sg13g2_decap_8
XFILLER_16_837 VPWR VGND sg13g2_decap_8
XFILLER_16_848 VPWR VGND sg13g2_fill_1
XFILLER_35_75 VPWR VGND sg13g2_fill_1
XFILLER_24_870 VPWR VGND sg13g2_fill_1
XFILLER_30_328 VPWR VGND sg13g2_fill_2
XFILLER_35_86 VPWR VGND sg13g2_decap_4
XFILLER_7_524 VPWR VGND sg13g2_decap_8
XFILLER_3_796 VPWR VGND sg13g2_decap_8
XFILLER_47_962 VPWR VGND sg13g2_decap_8
XFILLER_46_461 VPWR VGND sg13g2_fill_2
XFILLER_46_450 VPWR VGND sg13g2_decap_8
XFILLER_46_494 VPWR VGND sg13g2_fill_1
XFILLER_46_483 VPWR VGND sg13g2_fill_2
XFILLER_19_686 VPWR VGND sg13g2_decap_8
XFILLER_19_697 VPWR VGND sg13g2_fill_2
X_6067__213 VPWR VGND net213 sg13g2_tiehi
XFILLER_34_612 VPWR VGND sg13g2_decap_8
X_4810_ s0.data_out\[15\]\[0\] s0.data_out\[16\]\[0\] net1152 _0535_ VPWR VGND sg13g2_mux2_1
X_5790_ VGND VPWR net1030 _1415_ _1416_ _1375_ sg13g2_a21oi_1
XFILLER_34_689 VPWR VGND sg13g2_fill_1
X_4741_ VGND VPWR _0381_ _0470_ _0471_ net1160 sg13g2_a21oi_1
X_4672_ net1306 net308 _0048_ VPWR VGND sg13g2_and2_1
X_3623_ _2032_ net977 net355 VPWR VGND sg13g2_nand2_1
XFILLER_30_895 VPWR VGND sg13g2_fill_1
X_3554_ net970 net1064 _1968_ VPWR VGND sg13g2_nor2b_1
X_3485_ VGND VPWR net994 _1905_ _1906_ _1877_ sg13g2_a21oi_1
X_5224_ VGND VPWR _0840_ _0909_ _0910_ net1117 sg13g2_a21oi_1
XFILLER_5_1007 VPWR VGND sg13g2_decap_8
X_5155_ _0847_ net1112 _0822_ _0848_ VPWR VGND sg13g2_a21o_1
X_4106_ _2465_ net944 VPWR VGND sg13g2_inv_2
XFILLER_38_940 VPWR VGND sg13g2_decap_8
X_5086_ _0785_ net477 net1131 VPWR VGND sg13g2_nand2b_1
X_4037_ _2404_ VPWR _2405_ VGND net1292 net392 sg13g2_o21ai_1
XFILLER_25_623 VPWR VGND sg13g2_decap_4
X_5988_ net26 VGND VPWR _0038_ s0.valid_out\[18\][0] clknet_leaf_33_clk sg13g2_dfrbpq_1
XFILLER_13_829 VPWR VGND sg13g2_fill_2
X_4939_ _0652_ net921 _0651_ VPWR VGND sg13g2_nand2_1
XFILLER_4_516 VPWR VGND sg13g2_fill_1
XFILLER_43_1024 VPWR VGND sg13g2_decap_4
XFILLER_0_733 VPWR VGND sg13g2_decap_8
XFILLER_48_759 VPWR VGND sg13g2_decap_8
XFILLER_29_962 VPWR VGND sg13g2_fill_2
XFILLER_29_995 VPWR VGND sg13g2_decap_8
XFILLER_44_976 VPWR VGND sg13g2_decap_8
XFILLER_31_626 VPWR VGND sg13g2_decap_8
XFILLER_30_125 VPWR VGND sg13g2_decap_8
XFILLER_30_136 VPWR VGND sg13g2_fill_2
XFILLER_31_648 VPWR VGND sg13g2_decap_8
XFILLER_31_659 VPWR VGND sg13g2_fill_1
XFILLER_30_158 VPWR VGND sg13g2_fill_1
XFILLER_12_884 VPWR VGND sg13g2_fill_1
XFILLER_7_68 VPWR VGND sg13g2_fill_1
X_3270_ net1220 _1706_ _0189_ VPWR VGND sg13g2_nor2_1
Xfanout1350 rst_n net1350 VPWR VGND sg13g2_buf_8
X_5911_ _1526_ net517 net1032 VPWR VGND sg13g2_nand2b_1
XFILLER_35_921 VPWR VGND sg13g2_fill_1
XFILLER_46_280 VPWR VGND sg13g2_fill_2
X_5842_ VGND VPWR _1464_ _1466_ _0162_ _1467_ sg13g2_a21oi_1
X_5984__31 VPWR VGND net31 sg13g2_tiehi
X_5773_ VGND VPWR _1318_ _1400_ _1401_ net1037 sg13g2_a21oi_1
X_4724_ _0456_ net456 net1165 VPWR VGND sg13g2_nand2b_1
X_4655_ VGND VPWR net1172 _0395_ _0396_ _0340_ sg13g2_a21oi_1
X_4586_ VPWR _0042_ _0331_ VGND sg13g2_inv_1
X_3606_ VGND VPWR net970 _2014_ _2015_ _1968_ sg13g2_a21oi_1
X_3537_ net970 s0.data_out\[3\]\[1\] _1953_ VPWR VGND sg13g2_and2_1
X_3468_ VGND VPWR net981 _1888_ _1889_ _1837_ sg13g2_a21oi_1
X_6187_ net83 VGND VPWR _0237_ s0.valid_out\[2\][0] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_5207_ s0.data_out\[12\]\[1\] s0.data_out\[13\]\[1\] net1120 _0895_ VPWR VGND sg13g2_mux2_1
X_3399_ _1828_ net915 _1827_ VPWR VGND sg13g2_nand2_1
X_5138_ s0.data_out\[14\]\[1\] s0.data_out\[13\]\[1\] net1119 _0831_ VPWR VGND sg13g2_mux2_1
XFILLER_45_718 VPWR VGND sg13g2_decap_8
XFILLER_44_206 VPWR VGND sg13g2_fill_1
X_5069_ net1220 _0765_ _0086_ VPWR VGND sg13g2_nor2_1
XFILLER_25_431 VPWR VGND sg13g2_fill_2
XFILLER_25_464 VPWR VGND sg13g2_fill_2
XFILLER_26_987 VPWR VGND sg13g2_decap_8
XFILLER_41_968 VPWR VGND sg13g2_decap_8
XFILLER_9_608 VPWR VGND sg13g2_fill_1
XFILLER_40_478 VPWR VGND sg13g2_decap_8
XFILLER_40_489 VPWR VGND sg13g2_fill_1
XFILLER_5_825 VPWR VGND sg13g2_decap_8
XFILLER_0_530 VPWR VGND sg13g2_decap_8
XFILLER_48_534 VPWR VGND sg13g2_decap_8
XFILLER_44_784 VPWR VGND sg13g2_decap_4
XFILLER_44_773 VPWR VGND sg13g2_fill_2
XFILLER_43_261 VPWR VGND sg13g2_fill_1
XFILLER_17_998 VPWR VGND sg13g2_decap_8
X_6064__216 VPWR VGND net216 sg13g2_tiehi
XFILLER_32_968 VPWR VGND sg13g2_decap_8
X_5981__34 VPWR VGND net34 sg13g2_tiehi
X_4440_ s0.data_out\[18\]\[2\] s0.data_out\[19\]\[2\] net1186 _2762_ VPWR VGND sg13g2_mux2_1
Xhold107 s0.data_out\[4\]\[3\] VPWR VGND net403 sg13g2_dlygate4sd3_1
XFILLER_7_195 VPWR VGND sg13g2_fill_2
Xhold118 s0.data_out\[19\]\[4\] VPWR VGND net414 sg13g2_dlygate4sd3_1
Xhold129 _2182_ VPWR VGND net425 sg13g2_dlygate4sd3_1
X_6110_ net167 VGND VPWR _0160_ s0.data_out\[9\]\[6\] clknet_leaf_18_clk sg13g2_dfrbpq_2
X_4371_ VGND VPWR net1178 _2698_ _2699_ _2636_ sg13g2_a21oi_1
X_3322_ VGND VPWR net996 net538 _1757_ _1756_ sg13g2_a21oi_1
X_6071__209 VPWR VGND net209 sg13g2_tiehi
X_3253_ _1592_ VPWR _1698_ VGND _1691_ _1693_ sg13g2_o21ai_1
X_6041_ net241 VGND VPWR _0091_ s0.data_out\[14\]\[4\] clknet_leaf_25_clk sg13g2_dfrbpq_2
X_3184_ VGND VPWR net1005 net539 _1632_ _1631_ sg13g2_a21oi_1
XFILLER_39_556 VPWR VGND sg13g2_fill_1
Xfanout1180 net1181 net1180 VPWR VGND sg13g2_buf_1
Xfanout1191 net1192 net1191 VPWR VGND sg13g2_buf_1
XFILLER_35_751 VPWR VGND sg13g2_decap_4
X_5825_ _1450_ VPWR _1451_ VGND net1033 _2490_ sg13g2_o21ai_1
XFILLER_22_434 VPWR VGND sg13g2_decap_4
XFILLER_23_957 VPWR VGND sg13g2_decap_8
XFILLER_10_618 VPWR VGND sg13g2_decap_8
X_5756_ s0.data_out\[8\]\[4\] s0.data_out\[9\]\[4\] net1042 _1386_ VPWR VGND sg13g2_mux2_1
XFILLER_22_489 VPWR VGND sg13g2_fill_1
X_5687_ s0.data_out\[10\]\[5\] s0.data_out\[9\]\[5\] net1043 _1332_ VPWR VGND sg13g2_mux2_1
X_4707_ VPWR _0053_ _0441_ VGND sg13g2_inv_1
X_4638_ _0379_ _0378_ net1262 _0363_ net1269 VPWR VGND sg13g2_a22oi_1
X_4569_ _0316_ VPWR _0317_ VGND _0312_ _0315_ sg13g2_o21ai_1
XFILLER_26_740 VPWR VGND sg13g2_decap_4
XFILLER_41_732 VPWR VGND sg13g2_fill_2
XFILLER_13_445 VPWR VGND sg13g2_decap_8
XFILLER_14_968 VPWR VGND sg13g2_decap_8
XFILLER_9_427 VPWR VGND sg13g2_decap_8
XFILLER_13_489 VPWR VGND sg13g2_fill_2
XFILLER_40_297 VPWR VGND sg13g2_fill_1
XFILLER_5_644 VPWR VGND sg13g2_decap_8
XFILLER_1_872 VPWR VGND sg13g2_decap_8
XFILLER_49_821 VPWR VGND sg13g2_decap_8
XFILLER_0_393 VPWR VGND sg13g2_decap_8
XFILLER_49_898 VPWR VGND sg13g2_decap_8
XFILLER_48_397 VPWR VGND sg13g2_fill_2
X_3940_ _2317_ VPWR _2318_ VGND _2313_ _2316_ sg13g2_o21ai_1
XFILLER_32_721 VPWR VGND sg13g2_decap_8
X_3871_ _2256_ net956 net590 VPWR VGND sg13g2_nand2_1
XFILLER_20_905 VPWR VGND sg13g2_decap_8
XFILLER_31_242 VPWR VGND sg13g2_fill_2
XFILLER_31_264 VPWR VGND sg13g2_decap_8
X_5610_ s0.data_out\[9\]\[3\] s0.data_out\[10\]\[3\] net1087 _1260_ VPWR VGND sg13g2_mux2_1
XFILLER_9_950 VPWR VGND sg13g2_decap_8
X_5541_ VPWR VGND net1266 _1194_ _1197_ net1270 _1198_ _1184_ sg13g2_a221oi_1
X_5472_ net1335 VPWR _1136_ VGND net939 _1135_ sg13g2_o21ai_1
X_4423_ net1290 _2742_ _0026_ VPWR VGND sg13g2_and2_1
X_4354_ VGND VPWR _2591_ _2682_ _2683_ net1194 sg13g2_a21oi_1
X_3305_ net992 s0.data_out\[5\]\[4\] _1742_ VPWR VGND sg13g2_and2_1
X_4285_ net1196 VPWR _2623_ VGND net1225 net1182 sg13g2_o21ai_1
X_6024_ net259 VGND VPWR _0074_ s0.valid_out\[15\][0] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_3236_ _1678_ _1679_ _1680_ _1681_ VPWR VGND sg13g2_nor3_1
X_3167_ net1002 net1062 _1617_ VPWR VGND sg13g2_nor2b_1
XFILLER_35_581 VPWR VGND sg13g2_decap_8
X_5808_ VGND VPWR _1434_ _1417_ net1213 sg13g2_or2_1
X_5739_ VPWR _0155_ _1371_ VGND sg13g2_inv_1
XFILLER_2_636 VPWR VGND sg13g2_decap_8
Xfanout951 s0.shift_out\[1\][0] net951 VPWR VGND sg13g2_buf_8
XFILLER_38_20 VPWR VGND sg13g2_fill_2
XFILLER_1_168 VPWR VGND sg13g2_fill_1
Xfanout940 net941 net940 VPWR VGND sg13g2_buf_2
Xfanout962 net964 net962 VPWR VGND sg13g2_buf_8
Xfanout995 net996 net995 VPWR VGND sg13g2_buf_8
Xfanout984 net985 net984 VPWR VGND sg13g2_buf_8
Xfanout973 net975 net973 VPWR VGND sg13g2_buf_8
XFILLER_38_42 VPWR VGND sg13g2_fill_1
XFILLER_46_824 VPWR VGND sg13g2_decap_8
XFILLER_18_526 VPWR VGND sg13g2_decap_8
XFILLER_45_345 VPWR VGND sg13g2_decap_8
XFILLER_18_537 VPWR VGND sg13g2_decap_8
XFILLER_13_242 VPWR VGND sg13g2_decap_8
XFILLER_14_765 VPWR VGND sg13g2_decap_4
XFILLER_13_253 VPWR VGND sg13g2_fill_1
X_6061__219 VPWR VGND net219 sg13g2_tiehi
XFILLER_10_982 VPWR VGND sg13g2_decap_8
Xclkload16 VPWR clkload16/Y clknet_leaf_20_clk VGND sg13g2_inv_1
XFILLER_6_975 VPWR VGND sg13g2_decap_8
X_4070_ VPWR VGND _2429_ _2430_ _2428_ net1211 _2431_ _2408_ sg13g2_a221oi_1
XFILLER_49_695 VPWR VGND sg13g2_decap_8
X_4972_ net1126 s0.data_out\[14\]\[4\] _0681_ VPWR VGND sg13g2_and2_1
X_3923_ _2299_ _2302_ net1293 _2303_ VPWR VGND sg13g2_nand3_1
XFILLER_20_702 VPWR VGND sg13g2_decap_4
X_3854_ _2184_ _2238_ _2239_ VPWR VGND sg13g2_and2_1
XFILLER_32_562 VPWR VGND sg13g2_fill_1
XFILLER_20_746 VPWR VGND sg13g2_fill_1
XFILLER_9_780 VPWR VGND sg13g2_decap_4
X_3785_ net949 s0.data_out\[1\]\[0\] _2178_ VPWR VGND sg13g2_and2_1
X_5524_ _1181_ net1084 net506 VPWR VGND sg13g2_nand2_1
X_5455_ _1121_ VPWR _1122_ VGND net1080 _1115_ sg13g2_o21ai_1
X_4406_ net1214 _2723_ _2729_ _2734_ VPWR VGND sg13g2_or3_1
X_5386_ VGND VPWR _0965_ _1055_ _1056_ net1105 sg13g2_a21oi_1
XFILLER_8_1027 VPWR VGND sg13g2_fill_2
X_4337_ s0.data_out\[19\]\[5\] s0.data_out\[20\]\[5\] net1200 _2668_ VPWR VGND sg13g2_mux2_1
X_4268_ _2607_ net1196 _2550_ _2608_ VPWR VGND sg13g2_a21o_1
X_6007_ net278 VGND VPWR _0057_ s0.data_out\[17\]\[6\] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_3219_ VPWR VGND _1662_ _1663_ _1658_ net1212 _1664_ _1653_ sg13g2_a221oi_1
XFILLER_28_802 VPWR VGND sg13g2_fill_1
X_4199_ net1195 net1057 _2543_ VPWR VGND sg13g2_nor2b_1
XFILLER_28_835 VPWR VGND sg13g2_fill_1
XFILLER_43_849 VPWR VGND sg13g2_decap_8
XFILLER_27_389 VPWR VGND sg13g2_fill_2
XFILLER_11_713 VPWR VGND sg13g2_fill_2
XFILLER_24_66 VPWR VGND sg13g2_decap_8
XFILLER_10_212 VPWR VGND sg13g2_decap_8
XFILLER_10_223 VPWR VGND sg13g2_fill_2
XFILLER_11_768 VPWR VGND sg13g2_fill_2
XFILLER_6_227 VPWR VGND sg13g2_decap_8
XFILLER_3_901 VPWR VGND sg13g2_decap_8
XFILLER_3_978 VPWR VGND sg13g2_decap_8
XFILLER_2_477 VPWR VGND sg13g2_decap_4
XFILLER_2_488 VPWR VGND sg13g2_fill_2
Xhold290 s0.data_out\[19\]\[5\] VPWR VGND net586 sg13g2_dlygate4sd3_1
Xheichips25_top_sorter_19 VPWR VGND uio_out[4] sg13g2_tielo
XFILLER_19_846 VPWR VGND sg13g2_fill_1
XFILLER_34_805 VPWR VGND sg13g2_decap_4
XFILLER_46_698 VPWR VGND sg13g2_decap_8
X_6106__171 VPWR VGND net171 sg13g2_tiehi
X_3570_ net972 net1054 _1982_ VPWR VGND sg13g2_nor2b_1
XFILLER_6_783 VPWR VGND sg13g2_fill_2
X_5240_ VGND VPWR _0862_ _0923_ _0924_ net1117 sg13g2_a21oi_1
XFILLER_39_2 VPWR VGND sg13g2_fill_1
X_5171_ _0863_ net1114 _0808_ _0864_ VPWR VGND sg13g2_a21o_1
X_4122_ VPWR _2481_ s0.data_out\[21\]\[1\] VGND sg13g2_inv_1
X_4053_ net1294 net344 _2417_ VPWR VGND sg13g2_nor2_1
XFILLER_28_109 VPWR VGND sg13g2_fill_1
XFILLER_49_492 VPWR VGND sg13g2_decap_8
X_6113__164 VPWR VGND net164 sg13g2_tiehi
XFILLER_36_175 VPWR VGND sg13g2_fill_2
XFILLER_36_197 VPWR VGND sg13g2_fill_1
X_4955_ _0666_ net921 _0665_ VPWR VGND sg13g2_nand2_1
X_3906_ _2289_ _2286_ _2288_ VPWR VGND sg13g2_nand2_1
X_4886_ VPWR VGND _0602_ _0598_ _0597_ net1213 _0603_ _0593_ sg13g2_a221oi_1
X_3837_ _2223_ VPWR _2224_ VGND _2219_ _2222_ sg13g2_o21ai_1
X_3768_ VGND VPWR _2165_ net1210 net311 sg13g2_or2_1
XFILLER_20_598 VPWR VGND sg13g2_fill_1
X_5507_ VPWR _0128_ _1166_ VGND sg13g2_inv_1
X_3699_ VGND VPWR net963 net349 _2099_ _2098_ sg13g2_a21oi_1
XFILLER_10_13 VPWR VGND sg13g2_fill_1
X_5438_ _1099_ VPWR _1107_ VGND net1265 _1081_ sg13g2_o21ai_1
Xfanout1009 net1011 net1009 VPWR VGND sg13g2_buf_8
XFILLER_0_915 VPWR VGND sg13g2_decap_8
X_5369_ _1041_ s0.data_out\[11\]\[5\] net1110 VPWR VGND sg13g2_nand2b_1
XFILLER_47_407 VPWR VGND sg13g2_decap_8
XFILLER_19_99 VPWR VGND sg13g2_decap_8
XFILLER_28_676 VPWR VGND sg13g2_fill_1
XFILLER_42_101 VPWR VGND sg13g2_fill_2
XFILLER_3_775 VPWR VGND sg13g2_decap_8
XFILLER_47_941 VPWR VGND sg13g2_decap_8
XFILLER_19_643 VPWR VGND sg13g2_decap_8
XFILLER_20_1025 VPWR VGND sg13g2_decap_4
XFILLER_34_657 VPWR VGND sg13g2_fill_1
X_4740_ _0470_ s0.data_out\[16\]\[7\] net1164 VPWR VGND sg13g2_nand2b_1
XFILLER_14_392 VPWR VGND sg13g2_decap_8
X_4671_ VGND VPWR _0406_ _0410_ _0047_ _0411_ sg13g2_a21oi_1
XFILLER_30_874 VPWR VGND sg13g2_fill_1
X_3622_ _2031_ _2028_ _2029_ _2030_ VPWR VGND sg13g2_and3_1
X_3553_ net970 s0.data_out\[3\]\[3\] _1967_ VPWR VGND sg13g2_and2_1
X_3484_ _1904_ net984 _1878_ _1905_ VPWR VGND sg13g2_a21o_1
XFILLER_44_0 VPWR VGND sg13g2_decap_8
X_5223_ _0909_ net472 net1121 VPWR VGND sg13g2_nand2b_1
X_5154_ s0.data_out\[14\]\[7\] s0.data_out\[13\]\[7\] net1119 _0847_ VPWR VGND sg13g2_mux2_1
X_4105_ _2464_ net1138 VPWR VGND sg13g2_inv_2
XFILLER_29_418 VPWR VGND sg13g2_fill_2
X_5085_ VPWR _0088_ _0784_ VGND sg13g2_inv_1
X_4036_ net1292 VPWR _2404_ VGND _2402_ _2403_ sg13g2_o21ai_1
XFILLER_38_996 VPWR VGND sg13g2_decap_8
XFILLER_24_112 VPWR VGND sg13g2_decap_4
X_5987_ net28 VGND VPWR net407 s0.was_valid_out\[18\][0] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_25_679 VPWR VGND sg13g2_decap_4
X_4938_ s0.data_out\[14\]\[0\] s0.data_out\[15\]\[0\] net1142 _0651_ VPWR VGND sg13g2_mux2_1
XFILLER_33_690 VPWR VGND sg13g2_fill_1
X_4869_ VGND VPWR net1135 net554 _0587_ _0586_ sg13g2_a21oi_1
XFILLER_21_852 VPWR VGND sg13g2_fill_1
XFILLER_21_56 VPWR VGND sg13g2_fill_2
XFILLER_0_712 VPWR VGND sg13g2_decap_8
XFILLER_43_1003 VPWR VGND sg13g2_decap_8
XFILLER_0_789 VPWR VGND sg13g2_decap_8
XFILLER_48_738 VPWR VGND sg13g2_decap_8
XFILLER_29_930 VPWR VGND sg13g2_fill_1
XFILLER_29_974 VPWR VGND sg13g2_decap_8
XFILLER_44_955 VPWR VGND sg13g2_decap_8
XFILLER_15_134 VPWR VGND sg13g2_decap_8
XFILLER_12_863 VPWR VGND sg13g2_fill_1
XFILLER_7_58 VPWR VGND sg13g2_fill_1
X_6103__174 VPWR VGND net174 sg13g2_tiehi
XFILLER_3_550 VPWR VGND sg13g2_decap_8
XFILLER_39_705 VPWR VGND sg13g2_fill_2
Xfanout1340 net1341 net1340 VPWR VGND sg13g2_buf_8
XFILLER_16_4 VPWR VGND sg13g2_fill_2
X_5910_ VPWR _0172_ _1525_ VGND sg13g2_inv_1
X_6110__167 VPWR VGND net167 sg13g2_tiehi
X_5841_ VGND VPWR _1467_ net1210 net314 sg13g2_or2_1
XFILLER_35_999 VPWR VGND sg13g2_decap_8
X_5772_ _1400_ s0.data_out\[8\]\[6\] net1042 VPWR VGND sg13g2_nand2b_1
XFILLER_22_638 VPWR VGND sg13g2_fill_1
X_4723_ VPWR _0055_ _0455_ VGND sg13g2_inv_1
X_4654_ _0394_ net1159 _0341_ _0395_ VPWR VGND sg13g2_a21o_1
X_4585_ _0330_ VPWR _0331_ VGND net1301 net478 sg13g2_o21ai_1
X_3605_ s0.data_out\[4\]\[3\] s0.data_out\[3\]\[3\] net979 _2014_ VPWR VGND sg13g2_mux2_1
X_3536_ _1952_ net914 _1951_ VPWR VGND sg13g2_nand2_1
XFILLER_27_1009 VPWR VGND sg13g2_decap_8
X_5206_ VPWR _0099_ _0894_ VGND sg13g2_inv_1
X_3467_ s0.data_out\[5\]\[1\] s0.data_out\[4\]\[1\] net987 _1888_ VPWR VGND sg13g2_mux2_1
X_6186_ net85 VGND VPWR _0236_ s0.was_valid_out\[2\][0] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_3398_ s0.data_out\[4\]\[0\] s0.data_out\[5\]\[0\] net997 _1827_ VPWR VGND sg13g2_mux2_1
X_5137_ net1270 _0829_ _0830_ VPWR VGND sg13g2_nor2_1
X_5068_ VGND VPWR _0766_ _0769_ _0085_ _0770_ sg13g2_a21oi_1
XFILLER_29_259 VPWR VGND sg13g2_decap_8
X_4019_ _2387_ net1247 _2392_ VPWR VGND sg13g2_xor2_1
XFILLER_41_947 VPWR VGND sg13g2_decap_8
X_5990__24 VPWR VGND net24 sg13g2_tiehi
XFILLER_12_148 VPWR VGND sg13g2_fill_1
XFILLER_21_671 VPWR VGND sg13g2_fill_1
XFILLER_4_314 VPWR VGND sg13g2_fill_2
XFILLER_10_1024 VPWR VGND sg13g2_decap_4
XFILLER_4_347 VPWR VGND sg13g2_fill_1
X_6057__224 VPWR VGND net224 sg13g2_tiehi
XFILLER_48_513 VPWR VGND sg13g2_decap_8
XFILLER_0_586 VPWR VGND sg13g2_decap_8
XFILLER_17_900 VPWR VGND sg13g2_fill_2
XFILLER_28_281 VPWR VGND sg13g2_fill_1
XFILLER_44_752 VPWR VGND sg13g2_decap_8
XFILLER_17_977 VPWR VGND sg13g2_decap_8
XFILLER_40_980 VPWR VGND sg13g2_decap_8
Xhold108 s0.data_out\[10\]\[0\] VPWR VGND net404 sg13g2_dlygate4sd3_1
X_4370_ s0.data_out\[20\]\[0\] s0.data_out\[19\]\[0\] net1186 _2698_ VPWR VGND sg13g2_mux2_1
Xhold119 s0.data_out\[5\]\[3\] VPWR VGND net415 sg13g2_dlygate4sd3_1
X_3321_ net996 net1051 _1756_ VPWR VGND sg13g2_nor2b_1
XFILLER_3_380 VPWR VGND sg13g2_decap_8
X_6040_ net242 VGND VPWR _0090_ s0.data_out\[14\]\[3\] clknet_leaf_29_clk sg13g2_dfrbpq_2
X_3252_ _1677_ _1678_ _1697_ VPWR VGND sg13g2_nor2_1
X_3183_ net1005 net1055 _1631_ VPWR VGND sg13g2_nor2b_1
Xfanout1192 net1194 net1192 VPWR VGND sg13g2_buf_1
Xfanout1181 net1185 net1181 VPWR VGND sg13g2_buf_8
Xfanout1170 net1172 net1170 VPWR VGND sg13g2_buf_8
XFILLER_26_218 VPWR VGND sg13g2_fill_2
X_5824_ _1450_ net1033 net482 VPWR VGND sg13g2_nand2_1
XFILLER_34_284 VPWR VGND sg13g2_fill_2
X_5755_ VPWR _0157_ _1385_ VGND sg13g2_inv_1
X_4706_ _0440_ VPWR _0441_ VGND _0436_ _0439_ sg13g2_o21ai_1
X_5686_ _1268_ _1330_ net1257 _1331_ VPWR VGND sg13g2_nand3_1
X_4637_ _0326_ _0377_ _0378_ VPWR VGND sg13g2_and2_1
X_4568_ _0316_ net1219 _2484_ VPWR VGND sg13g2_nand2_1
X_3519_ net353 _1937_ _1938_ VPWR VGND sg13g2_nor2_1
X_4499_ VGND VPWR net1167 _2814_ _2815_ _2751_ sg13g2_a21oi_1
X_6169_ net103 VGND VPWR _0219_ s0.data_out\[4\]\[5\] clknet_leaf_12_clk sg13g2_dfrbpq_2
XFILLER_18_708 VPWR VGND sg13g2_decap_8
XFILLER_17_218 VPWR VGND sg13g2_fill_1
XFILLER_18_719 VPWR VGND sg13g2_fill_1
XFILLER_25_240 VPWR VGND sg13g2_fill_1
XFILLER_14_925 VPWR VGND sg13g2_fill_1
X_6208__260 VPWR VGND net260 sg13g2_tiehi
XFILLER_40_243 VPWR VGND sg13g2_decap_8
XFILLER_40_221 VPWR VGND sg13g2_fill_2
XFILLER_43_76 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_20_clk clknet_3_7__leaf_clk clknet_leaf_20_clk VPWR VGND sg13g2_buf_8
XFILLER_4_188 VPWR VGND sg13g2_fill_2
XFILLER_49_800 VPWR VGND sg13g2_decap_8
XFILLER_1_851 VPWR VGND sg13g2_decap_8
X_6070__210 VPWR VGND net210 sg13g2_tiehi
XFILLER_49_877 VPWR VGND sg13g2_decap_8
XFILLER_17_774 VPWR VGND sg13g2_decap_4
XFILLER_17_796 VPWR VGND sg13g2_fill_2
X_3870_ VGND VPWR net964 _2254_ _2255_ _2226_ sg13g2_a21oi_1
XFILLER_17_1019 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_11_clk clknet_3_3__leaf_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
XFILLER_13_991 VPWR VGND sg13g2_decap_8
X_5540_ VGND VPWR net1095 _1196_ _1197_ _1147_ sg13g2_a21oi_1
XFILLER_31_298 VPWR VGND sg13g2_decap_4
X_5471_ VGND VPWR net1077 net418 _1135_ _1134_ sg13g2_a21oi_1
X_4422_ VGND VPWR _2447_ _2742_ _0025_ _2747_ sg13g2_a21oi_1
X_4353_ _2682_ s0.data_out\[19\]\[7\] net1199 VPWR VGND sg13g2_nand2b_1
X_4284_ net1285 net301 _0012_ VPWR VGND sg13g2_and2_1
X_3304_ _1741_ net916 _1740_ VPWR VGND sg13g2_nand2_1
X_6023_ net261 VGND VPWR net382 s0.was_valid_out\[15\][0] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_3235_ net1264 _1667_ _1680_ VPWR VGND sg13g2_nor2_1
XFILLER_39_332 VPWR VGND sg13g2_decap_4
XFILLER_27_505 VPWR VGND sg13g2_fill_2
X_3166_ VGND VPWR _1545_ _1615_ _1616_ net1012 sg13g2_a21oi_1
XFILLER_39_398 VPWR VGND sg13g2_fill_1
X_3999_ s0.data_out\[1\]\[6\] s0.data_out\[0\]\[6\] net947 _2372_ VPWR VGND sg13g2_mux2_1
XFILLER_22_254 VPWR VGND sg13g2_fill_1
X_5807_ _1433_ net1266 _1432_ VPWR VGND sg13g2_nand2_1
XFILLER_10_438 VPWR VGND sg13g2_decap_4
X_5738_ _1370_ VPWR _1371_ VGND net1340 net405 sg13g2_o21ai_1
X_5669_ _1314_ net1043 net565 VPWR VGND sg13g2_nand2_1
XFILLER_2_615 VPWR VGND sg13g2_decap_8
X_6054__227 VPWR VGND net227 sg13g2_tiehi
Xfanout952 net954 net952 VPWR VGND sg13g2_buf_8
Xfanout930 _2458_ net930 VPWR VGND sg13g2_buf_8
Xfanout941 net942 net941 VPWR VGND sg13g2_buf_2
Xfanout963 net964 net963 VPWR VGND sg13g2_buf_8
Xfanout985 net986 net985 VPWR VGND sg13g2_buf_8
Xfanout974 net975 net974 VPWR VGND sg13g2_buf_1
XFILLER_46_803 VPWR VGND sg13g2_decap_8
Xfanout996 s0.shift_out\[5\][0] net996 VPWR VGND sg13g2_buf_8
XFILLER_45_313 VPWR VGND sg13g2_fill_1
XFILLER_10_961 VPWR VGND sg13g2_decap_8
Xclkload17 VPWR clkload17/Y clknet_leaf_21_clk VGND sg13g2_inv_1
XFILLER_6_954 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_49_674 VPWR VGND sg13g2_decap_8
XFILLER_37_814 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_0_clk clknet_3_0__leaf_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
XFILLER_36_379 VPWR VGND sg13g2_decap_4
X_4971_ _0680_ _2464_ _0679_ VPWR VGND sg13g2_nand2_1
XFILLER_17_582 VPWR VGND sg13g2_decap_8
X_3922_ net951 VPWR _2302_ VGND _2300_ _2301_ sg13g2_o21ai_1
XFILLER_32_530 VPWR VGND sg13g2_fill_2
X_3853_ _2238_ net961 _2237_ VPWR VGND sg13g2_nand2b_1
X_3784_ _2177_ net930 _2176_ VPWR VGND sg13g2_nand2_1
XFILLER_30_1016 VPWR VGND sg13g2_decap_8
X_5523_ VPWR _0130_ _1180_ VGND sg13g2_inv_1
XFILLER_30_1027 VPWR VGND sg13g2_fill_2
X_5454_ net939 VPWR _1121_ VGND net379 net1097 sg13g2_o21ai_1
X_4405_ _2720_ _2728_ _2731_ _2732_ _2733_ VPWR VGND sg13g2_and4_1
X_5385_ _1055_ net540 net1110 VPWR VGND sg13g2_nand2b_1
XFILLER_5_80 VPWR VGND sg13g2_decap_4
XFILLER_8_1006 VPWR VGND sg13g2_decap_8
X_4336_ VPWR _0019_ _2667_ VGND sg13g2_inv_1
X_4267_ s0.data_out\[21\]\[5\] s0.data_out\[20\]\[5\] net1200 _2607_ VPWR VGND sg13g2_mux2_1
X_4198_ net1196 s0.data_out\[20\]\[4\] _2542_ VPWR VGND sg13g2_and2_1
X_6006_ net279 VGND VPWR _0056_ s0.data_out\[17\]\[5\] clknet_leaf_32_clk sg13g2_dfrbpq_2
XFILLER_27_302 VPWR VGND sg13g2_fill_2
X_3218_ VGND VPWR _1602_ _1657_ _1663_ net1278 sg13g2_a21oi_1
XFILLER_39_184 VPWR VGND sg13g2_fill_2
X_3149_ s0.data_out\[6\]\[1\] s0.data_out\[7\]\[1\] net1019 _1601_ VPWR VGND sg13g2_mux2_1
XFILLER_27_346 VPWR VGND sg13g2_fill_2
XFILLER_42_349 VPWR VGND sg13g2_decap_8
X_6060__220 VPWR VGND net220 sg13g2_tiehi
XFILLER_40_88 VPWR VGND sg13g2_decap_8
Xhold280 s0.data_out\[3\]\[6\] VPWR VGND net576 sg13g2_dlygate4sd3_1
XFILLER_3_957 VPWR VGND sg13g2_decap_8
XFILLER_2_445 VPWR VGND sg13g2_decap_8
XFILLER_49_42 VPWR VGND sg13g2_decap_8
Xhold291 s0.data_out\[8\]\[6\] VPWR VGND net587 sg13g2_dlygate4sd3_1
XFILLER_46_677 VPWR VGND sg13g2_decap_8
XFILLER_14_552 VPWR VGND sg13g2_fill_2
XFILLER_42_894 VPWR VGND sg13g2_decap_8
X_6217__123 VPWR VGND net123 sg13g2_tiehi
X_5170_ s0.data_out\[14\]\[5\] s0.data_out\[13\]\[5\] net1120 _0863_ VPWR VGND sg13g2_mux2_1
X_4121_ _2480_ net1268 VPWR VGND sg13g2_inv_2
X_4052_ VPWR _0266_ _2416_ VGND sg13g2_inv_1
XFILLER_49_471 VPWR VGND sg13g2_decap_8
XFILLER_37_666 VPWR VGND sg13g2_fill_1
X_4954_ s0.data_out\[14\]\[2\] s0.data_out\[15\]\[2\] net1142 _0665_ VPWR VGND sg13g2_mux2_1
X_3905_ net929 VPWR _2288_ VGND s0.was_valid_out\[0\][0] net956 sg13g2_o21ai_1
X_4885_ net1282 _0601_ _0602_ VPWR VGND sg13g2_nor2b_1
X_3836_ VGND VPWR _2223_ net491 net1299 sg13g2_or2_1
X_3767_ _2055_ _2162_ _2163_ _2164_ VPWR VGND sg13g2_nor3_1
X_5506_ _1165_ VPWR _1166_ VGND _1161_ _1164_ sg13g2_o21ai_1
X_3698_ net963 net1054 _2098_ VPWR VGND sg13g2_nor2b_1
XFILLER_10_69 VPWR VGND sg13g2_decap_8
X_5437_ VGND VPWR _1106_ _1098_ net1256 sg13g2_or2_1
X_5368_ VPWR _0115_ _1040_ VGND sg13g2_inv_1
X_4319_ _2652_ VPWR _2653_ VGND _2648_ _2651_ sg13g2_o21ai_1
X_5299_ VGND VPWR net1102 _0979_ _0980_ _0919_ sg13g2_a21oi_1
XFILLER_28_611 VPWR VGND sg13g2_fill_1
XFILLER_15_327 VPWR VGND sg13g2_fill_2
XFILLER_27_187 VPWR VGND sg13g2_fill_1
XFILLER_11_500 VPWR VGND sg13g2_fill_2
XFILLER_11_577 VPWR VGND sg13g2_decap_8
XFILLER_11_588 VPWR VGND sg13g2_fill_1
X_5999__287 VPWR VGND net287 sg13g2_tiehi
XFILLER_3_754 VPWR VGND sg13g2_decap_8
XFILLER_2_253 VPWR VGND sg13g2_fill_1
XFILLER_2_286 VPWR VGND sg13g2_fill_1
XFILLER_47_920 VPWR VGND sg13g2_decap_8
XFILLER_19_633 VPWR VGND sg13g2_fill_1
XFILLER_20_1004 VPWR VGND sg13g2_decap_8
XFILLER_18_110 VPWR VGND sg13g2_decap_4
XFILLER_47_997 VPWR VGND sg13g2_decap_8
XFILLER_46_485 VPWR VGND sg13g2_fill_1
XFILLER_33_124 VPWR VGND sg13g2_fill_1
XFILLER_14_371 VPWR VGND sg13g2_fill_2
X_4670_ VGND VPWR _0411_ net1210 net304 sg13g2_or2_1
X_3621_ VGND VPWR _2030_ _2023_ net1234 sg13g2_or2_1
X_3552_ _1966_ net914 _1965_ VPWR VGND sg13g2_nand2_1
XFILLER_6_581 VPWR VGND sg13g2_decap_4
X_3483_ s0.data_out\[5\]\[7\] s0.data_out\[4\]\[7\] net988 _1904_ VPWR VGND sg13g2_mux2_1
X_5222_ VPWR _0101_ _0908_ VGND sg13g2_inv_1
XFILLER_37_0 VPWR VGND sg13g2_decap_4
X_5153_ _0846_ net1121 net584 VPWR VGND sg13g2_nand2_1
X_4104_ VPWR _2463_ net1148 VGND sg13g2_inv_1
X_5084_ _0783_ VPWR _0784_ VGND _0779_ _0782_ sg13g2_o21ai_1
XFILLER_38_975 VPWR VGND sg13g2_decap_8
XFILLER_2_92 VPWR VGND sg13g2_fill_2
X_4035_ net1069 net940 _2403_ VPWR VGND sg13g2_nor2b_1
X_5986_ net29 VGND VPWR _0036_ s0.genblk1\[18\].modules.bubble clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_36_1022 VPWR VGND sg13g2_decap_8
X_4937_ net1220 _0645_ _0074_ VPWR VGND sg13g2_nor2_1
X_4868_ net1135 net1047 _0586_ VPWR VGND sg13g2_nor2b_1
X_3819_ net962 VPWR _2208_ VGND _2206_ _2207_ sg13g2_o21ai_1
XFILLER_21_886 VPWR VGND sg13g2_fill_2
X_4799_ net1228 net1143 _0526_ VPWR VGND sg13g2_nor2b_1
XFILLER_21_46 VPWR VGND sg13g2_decap_4
XFILLER_48_717 VPWR VGND sg13g2_decap_8
XFILLER_0_768 VPWR VGND sg13g2_decap_8
XFILLER_29_964 VPWR VGND sg13g2_fill_1
XFILLER_44_934 VPWR VGND sg13g2_decap_8
XFILLER_43_400 VPWR VGND sg13g2_decap_8
X_6219__97 VPWR VGND net97 sg13g2_tiehi
XFILLER_16_625 VPWR VGND sg13g2_decap_8
XFILLER_43_455 VPWR VGND sg13g2_decap_4
XFILLER_15_146 VPWR VGND sg13g2_decap_8
XFILLER_7_301 VPWR VGND sg13g2_fill_2
XFILLER_11_363 VPWR VGND sg13g2_decap_4
XFILLER_7_345 VPWR VGND sg13g2_decap_8
XFILLER_7_389 VPWR VGND sg13g2_fill_2
XFILLER_30_7 VPWR VGND sg13g2_fill_2
Xfanout1330 net1331 net1330 VPWR VGND sg13g2_buf_1
Xfanout1341 net1348 net1341 VPWR VGND sg13g2_buf_8
XFILLER_34_400 VPWR VGND sg13g2_fill_1
XFILLER_47_794 VPWR VGND sg13g2_decap_8
XFILLER_34_411 VPWR VGND sg13g2_fill_1
X_5840_ VPWR VGND _1465_ _1352_ _1449_ _1445_ _1466_ _1447_ sg13g2_a221oi_1
XFILLER_35_978 VPWR VGND sg13g2_decap_8
X_5771_ VPWR _0159_ _1399_ VGND sg13g2_inv_1
XFILLER_21_105 VPWR VGND sg13g2_fill_1
X_4722_ _0454_ VPWR _0455_ VGND net1306 net401 sg13g2_o21ai_1
X_4653_ s0.data_out\[18\]\[5\] s0.data_out\[17\]\[5\] net1166 _0394_ VPWR VGND sg13g2_mux2_1
X_4584_ _0326_ _0329_ net1301 _0330_ VPWR VGND sg13g2_nand3_1
X_3604_ _2013_ net976 net509 VPWR VGND sg13g2_nand2_1
X_3535_ s0.data_out\[3\]\[1\] s0.data_out\[4\]\[1\] net987 _1951_ VPWR VGND sg13g2_mux2_1
X_3466_ VGND VPWR _1887_ _1886_ net1271 sg13g2_or2_1
X_5205_ _0893_ VPWR _0894_ VGND net1333 net439 sg13g2_o21ai_1
X_6185_ net86 VGND VPWR _0235_ s0.genblk1\[2\].modules.bubble clknet_leaf_10_clk sg13g2_dfrbpq_1
X_3397_ net1219 _1821_ _0201_ VPWR VGND sg13g2_nor2_1
X_5136_ VGND VPWR net1127 _0828_ _0829_ _0786_ sg13g2_a21oi_1
X_5067_ net1321 VPWR _0770_ VGND net378 _0765_ sg13g2_o21ai_1
XFILLER_29_238 VPWR VGND sg13g2_decap_8
XFILLER_37_260 VPWR VGND sg13g2_decap_8
X_4018_ _2391_ net1254 _2382_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_794 VPWR VGND sg13g2_fill_1
XFILLER_25_433 VPWR VGND sg13g2_fill_1
XFILLER_26_967 VPWR VGND sg13g2_decap_4
XFILLER_41_926 VPWR VGND sg13g2_decap_8
XFILLER_16_68 VPWR VGND sg13g2_decap_8
XFILLER_25_444 VPWR VGND sg13g2_decap_4
XFILLER_25_466 VPWR VGND sg13g2_fill_1
XFILLER_12_105 VPWR VGND sg13g2_fill_1
XFILLER_12_116 VPWR VGND sg13g2_fill_2
X_5969_ net47 VGND VPWR _0019_ s0.data_out\[20\]\[4\] clknet_leaf_2_clk sg13g2_dfrbpq_2
XFILLER_21_661 VPWR VGND sg13g2_fill_2
XFILLER_20_182 VPWR VGND sg13g2_decap_8
XFILLER_10_1003 VPWR VGND sg13g2_decap_8
XFILLER_0_565 VPWR VGND sg13g2_decap_8
XFILLER_48_547 VPWR VGND sg13g2_decap_8
XFILLER_17_934 VPWR VGND sg13g2_fill_1
XFILLER_16_488 VPWR VGND sg13g2_fill_1
XFILLER_16_499 VPWR VGND sg13g2_decap_8
XFILLER_31_425 VPWR VGND sg13g2_fill_1
XFILLER_43_296 VPWR VGND sg13g2_fill_1
XFILLER_31_458 VPWR VGND sg13g2_fill_1
XFILLER_31_469 VPWR VGND sg13g2_fill_2
XFILLER_7_197 VPWR VGND sg13g2_fill_1
Xhold109 s0.data_out\[9\]\[1\] VPWR VGND net405 sg13g2_dlygate4sd3_1
X_3320_ VGND VPWR _1687_ _1754_ _1755_ net1004 sg13g2_a21oi_1
XFILLER_4_893 VPWR VGND sg13g2_decap_8
X_3251_ _1695_ VPWR _1696_ VGND _1664_ _1669_ sg13g2_o21ai_1
X_3182_ VGND VPWR _1569_ _1629_ _1630_ net1015 sg13g2_a21oi_1
XFILLER_39_503 VPWR VGND sg13g2_decap_8
Xfanout1160 net1161 net1160 VPWR VGND sg13g2_buf_8
Xfanout1171 net1172 net1171 VPWR VGND sg13g2_buf_8
Xfanout1182 net1183 net1182 VPWR VGND sg13g2_buf_8
Xfanout1193 net1194 net1193 VPWR VGND sg13g2_buf_8
XFILLER_35_775 VPWR VGND sg13g2_fill_2
X_5823_ _1446_ _1448_ _1449_ VPWR VGND sg13g2_nor2_1
XFILLER_34_263 VPWR VGND sg13g2_fill_1
X_5754_ _1384_ VPWR _1385_ VGND net1340 net400 sg13g2_o21ai_1
XFILLER_33_1025 VPWR VGND sg13g2_decap_4
X_4705_ VGND VPWR _0440_ net530 net1304 sg13g2_or2_1
XFILLER_30_491 VPWR VGND sg13g2_fill_1
XFILLER_31_992 VPWR VGND sg13g2_decap_8
X_5685_ _1330_ net1082 _1329_ VPWR VGND sg13g2_nand2b_1
X_4636_ _0377_ net1169 _0376_ VPWR VGND sg13g2_nand2b_1
XFILLER_2_819 VPWR VGND sg13g2_decap_8
X_4567_ net1301 VPWR _0315_ VGND net925 _0314_ sg13g2_o21ai_1
X_3518_ _1936_ VPWR _1937_ VGND net983 _1818_ sg13g2_o21ai_1
X_4498_ s0.data_out\[19\]\[0\] s0.data_out\[18\]\[0\] net1174 _2814_ VPWR VGND sg13g2_mux2_1
X_3449_ VGND VPWR net985 net511 _1872_ _1871_ sg13g2_a21oi_1
X_6168_ net104 VGND VPWR _0218_ s0.data_out\[4\]\[4\] clknet_leaf_14_clk sg13g2_dfrbpq_2
X_5119_ VGND VPWR _0733_ _0813_ _0814_ net1128 sg13g2_a21oi_1
X_6099_ net179 VGND VPWR _0149_ s0.data_new_delayed\[5\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_41_734 VPWR VGND sg13g2_fill_1
XFILLER_40_200 VPWR VGND sg13g2_decap_8
XFILLER_25_252 VPWR VGND sg13g2_fill_2
XFILLER_26_797 VPWR VGND sg13g2_decap_8
XFILLER_43_55 VPWR VGND sg13g2_decap_4
XFILLER_40_233 VPWR VGND sg13g2_fill_1
XFILLER_21_491 VPWR VGND sg13g2_decap_8
XFILLER_22_992 VPWR VGND sg13g2_decap_8
XFILLER_49_1010 VPWR VGND sg13g2_decap_8
XFILLER_4_145 VPWR VGND sg13g2_fill_2
XFILLER_4_134 VPWR VGND sg13g2_decap_8
X_6100__178 VPWR VGND net178 sg13g2_tiehi
XFILLER_4_27 VPWR VGND sg13g2_fill_2
XFILLER_1_830 VPWR VGND sg13g2_decap_8
XFILLER_0_362 VPWR VGND sg13g2_decap_8
XFILLER_0_373 VPWR VGND sg13g2_fill_2
XFILLER_49_856 VPWR VGND sg13g2_decap_8
XFILLER_36_539 VPWR VGND sg13g2_fill_1
XFILLER_1_1012 VPWR VGND sg13g2_decap_8
XFILLER_29_591 VPWR VGND sg13g2_fill_1
XFILLER_16_274 VPWR VGND sg13g2_fill_1
XFILLER_31_211 VPWR VGND sg13g2_fill_2
XFILLER_32_767 VPWR VGND sg13g2_fill_2
XFILLER_13_970 VPWR VGND sg13g2_decap_8
XFILLER_9_985 VPWR VGND sg13g2_decap_8
X_5470_ net1077 net1070 _1134_ VPWR VGND sg13g2_nor2b_1
XFILLER_8_484 VPWR VGND sg13g2_fill_2
X_4421_ net1290 VPWR _2747_ VGND _2744_ _2746_ sg13g2_o21ai_1
X_4352_ VPWR _0021_ _2681_ VGND sg13g2_inv_1
X_4283_ VGND VPWR _2616_ _2620_ _0011_ _2622_ sg13g2_a21oi_1
X_3303_ s0.data_out\[5\]\[4\] s0.data_out\[6\]\[4\] net1008 _1740_ VPWR VGND sg13g2_mux2_1
X_6022_ net262 VGND VPWR _0072_ s0.genblk1\[15\].modules.bubble clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
X_3234_ net1258 _1672_ _1679_ VPWR VGND sg13g2_nor2_1
X_3165_ _1615_ net454 net1019 VPWR VGND sg13g2_nand2b_1
XFILLER_42_509 VPWR VGND sg13g2_fill_2
XFILLER_35_561 VPWR VGND sg13g2_fill_2
XFILLER_11_907 VPWR VGND sg13g2_fill_2
X_6047__235 VPWR VGND net235 sg13g2_tiehi
X_3998_ VGND VPWR net954 _2370_ _2371_ _2341_ sg13g2_a21oi_1
XFILLER_10_417 VPWR VGND sg13g2_fill_1
X_5806_ _1380_ _1431_ _1432_ VPWR VGND sg13g2_and2_1
XFILLER_22_288 VPWR VGND sg13g2_decap_4
X_5737_ _1366_ _1369_ net1341 _1370_ VPWR VGND sg13g2_nand3_1
XFILLER_13_58 VPWR VGND sg13g2_fill_1
X_5668_ _1312_ VPWR _1313_ VGND _1306_ _1307_ sg13g2_o21ai_1
X_4619_ _0360_ net1164 net530 VPWR VGND sg13g2_nand2_1
X_5599_ _1247_ _1250_ net1341 _1251_ VPWR VGND sg13g2_nand3_1
XFILLER_49_119 VPWR VGND sg13g2_decap_8
Xfanout920 _2466_ net920 VPWR VGND sg13g2_buf_1
Xfanout942 net945 net942 VPWR VGND sg13g2_buf_8
XFILLER_1_159 VPWR VGND sg13g2_decap_8
Xfanout931 _2456_ net931 VPWR VGND sg13g2_buf_8
Xfanout964 s0.shift_out\[2\][0] net964 VPWR VGND sg13g2_buf_8
Xfanout953 net954 net953 VPWR VGND sg13g2_buf_8
Xfanout986 s0.shift_out\[4\][0] net986 VPWR VGND sg13g2_buf_8
Xfanout975 s0.shift_out\[3\][0] net975 VPWR VGND sg13g2_buf_8
Xfanout997 net999 net997 VPWR VGND sg13g2_buf_8
XFILLER_46_859 VPWR VGND sg13g2_decap_8
XFILLER_38_99 VPWR VGND sg13g2_fill_1
XFILLER_26_561 VPWR VGND sg13g2_decap_8
XFILLER_14_734 VPWR VGND sg13g2_decap_8
XFILLER_26_594 VPWR VGND sg13g2_fill_1
XFILLER_10_940 VPWR VGND sg13g2_decap_8
XFILLER_6_933 VPWR VGND sg13g2_decap_8
XFILLER_23_1013 VPWR VGND sg13g2_decap_8
XFILLER_49_653 VPWR VGND sg13g2_decap_8
XFILLER_48_130 VPWR VGND sg13g2_fill_2
XFILLER_0_192 VPWR VGND sg13g2_decap_8
XFILLER_24_509 VPWR VGND sg13g2_fill_1
XFILLER_17_561 VPWR VGND sg13g2_fill_2
X_4970_ s0.data_out\[14\]\[4\] s0.data_out\[15\]\[4\] net1143 _0679_ VPWR VGND sg13g2_mux2_1
X_3921_ net942 net1069 _2301_ VPWR VGND sg13g2_nor2b_1
X_3852_ VGND VPWR net949 _2236_ _2237_ _2186_ sg13g2_a21oi_1
X_3783_ s0.data_out\[1\]\[0\] s0.data_out\[2\]\[0\] net965 _2176_ VPWR VGND sg13g2_mux2_1
X_5522_ _1179_ VPWR _1180_ VGND _1175_ _1178_ sg13g2_o21ai_1
X_5453_ VGND VPWR _1120_ net1085 net379 sg13g2_or2_1
X_4404_ _2732_ net1254 _2723_ VPWR VGND sg13g2_xnor2_1
X_5384_ VPWR _0117_ _1054_ VGND sg13g2_inv_1
X_4335_ _2666_ VPWR _2667_ VGND net1289 net469 sg13g2_o21ai_1
X_4266_ _2606_ net1254 _2605_ VPWR VGND sg13g2_nand2_1
X_4197_ _0006_ _2537_ _2541_ _2478_ net1216 VPWR VGND sg13g2_a22oi_1
X_6005_ net280 VGND VPWR _0055_ s0.data_out\[17\]\[4\] clknet_leaf_4_clk sg13g2_dfrbpq_2
X_3217_ net1282 _1661_ _1662_ VPWR VGND sg13g2_nor2b_1
X_3148_ VPWR _0178_ _1600_ VGND sg13g2_inv_1
XFILLER_27_314 VPWR VGND sg13g2_fill_2
XFILLER_43_818 VPWR VGND sg13g2_decap_8
XFILLER_23_553 VPWR VGND sg13g2_fill_2
XFILLER_11_726 VPWR VGND sg13g2_decap_8
XFILLER_40_12 VPWR VGND sg13g2_decap_8
XFILLER_40_78 VPWR VGND sg13g2_fill_1
XFILLER_40_56 VPWR VGND sg13g2_decap_4
XFILLER_3_936 VPWR VGND sg13g2_decap_8
XFILLER_49_21 VPWR VGND sg13g2_decap_8
XFILLER_46_1013 VPWR VGND sg13g2_decap_8
Xhold270 _1413_ VPWR VGND net566 sg13g2_dlygate4sd3_1
XFILLER_6_4 VPWR VGND sg13g2_fill_2
Xhold281 s0.data_out\[14\]\[7\] VPWR VGND net577 sg13g2_dlygate4sd3_1
Xhold292 s0.data_out\[12\]\[6\] VPWR VGND net588 sg13g2_dlygate4sd3_1
XFILLER_49_98 VPWR VGND sg13g2_decap_8
XFILLER_19_837 VPWR VGND sg13g2_decap_8
XFILLER_46_656 VPWR VGND sg13g2_decap_8
XFILLER_18_336 VPWR VGND sg13g2_decap_4
XFILLER_45_166 VPWR VGND sg13g2_fill_2
XFILLER_27_892 VPWR VGND sg13g2_fill_2
XFILLER_42_873 VPWR VGND sg13g2_decap_8
XFILLER_14_586 VPWR VGND sg13g2_fill_2
XFILLER_5_262 VPWR VGND sg13g2_decap_8
XFILLER_5_295 VPWR VGND sg13g2_fill_2
X_6037__245 VPWR VGND net245 sg13g2_tiehi
X_4120_ VPWR _2479_ s0.data_out\[21\]\[2\] VGND sg13g2_inv_1
XFILLER_2_980 VPWR VGND sg13g2_decap_8
XFILLER_49_450 VPWR VGND sg13g2_decap_8
XFILLER_1_490 VPWR VGND sg13g2_decap_4
X_4051_ VGND VPWR net1218 net374 _2416_ _2415_ sg13g2_a21oi_1
XFILLER_37_645 VPWR VGND sg13g2_fill_2
XFILLER_36_133 VPWR VGND sg13g2_decap_4
XFILLER_18_881 VPWR VGND sg13g2_decap_8
X_4953_ VPWR _0076_ _0664_ VGND sg13g2_inv_1
XFILLER_24_328 VPWR VGND sg13g2_decap_4
XFILLER_33_840 VPWR VGND sg13g2_fill_1
X_3904_ net943 _2283_ _2287_ VPWR VGND sg13g2_nor2_1
X_6044__238 VPWR VGND net238 sg13g2_tiehi
X_4884_ _0536_ VPWR _0601_ VGND net922 _0600_ sg13g2_o21ai_1
XFILLER_32_383 VPWR VGND sg13g2_fill_2
X_3835_ net1299 VPWR _2222_ VGND _2458_ _2221_ sg13g2_o21ai_1
X_3766_ _2144_ _2146_ _2163_ VPWR VGND sg13g2_nor2b_1
X_5505_ VGND VPWR _1165_ net541 net1336 sg13g2_or2_1
X_3697_ VGND VPWR _2032_ _2096_ _2097_ net973 sg13g2_a21oi_1
X_5436_ VGND VPWR _1105_ _1103_ net1251 sg13g2_or2_1
X_5367_ _1039_ VPWR _1040_ VGND net331 _1038_ sg13g2_o21ai_1
X_4318_ VGND VPWR _2652_ net490 net1285 sg13g2_or2_1
X_5298_ s0.data_out\[13\]\[4\] s0.data_out\[12\]\[4\] net1108 _0979_ VPWR VGND sg13g2_mux2_1
X_4249_ _2588_ VPWR _2589_ VGND net1211 _2573_ sg13g2_o21ai_1
XFILLER_28_645 VPWR VGND sg13g2_decap_8
XFILLER_28_667 VPWR VGND sg13g2_decap_8
XFILLER_43_604 VPWR VGND sg13g2_decap_4
XFILLER_23_372 VPWR VGND sg13g2_decap_4
XFILLER_13_1012 VPWR VGND sg13g2_decap_8
XFILLER_3_733 VPWR VGND sg13g2_decap_8
XFILLER_2_243 VPWR VGND sg13g2_fill_1
XFILLER_47_976 VPWR VGND sg13g2_decap_8
XFILLER_21_309 VPWR VGND sg13g2_decap_8
X_3620_ VGND VPWR _2029_ _2027_ net1241 sg13g2_or2_1
X_3551_ s0.data_out\[3\]\[3\] s0.data_out\[4\]\[3\] net987 _1965_ VPWR VGND sg13g2_mux2_1
X_3482_ _1903_ net988 net535 VPWR VGND sg13g2_nand2_1
X_5221_ _0907_ VPWR _0908_ VGND net1332 net477 sg13g2_o21ai_1
X_5152_ VPWR VGND net1265 _0839_ _0844_ net1270 _0845_ _0829_ sg13g2_a221oi_1
X_4103_ _2462_ net1160 VPWR VGND sg13g2_inv_2
X_5083_ VGND VPWR _0783_ net564 net1320 sg13g2_or2_1
X_6050__231 VPWR VGND net231 sg13g2_tiehi
XFILLER_38_954 VPWR VGND sg13g2_decap_8
X_4034_ VGND VPWR net946 net392 _2402_ net940 sg13g2_a21oi_1
XFILLER_25_648 VPWR VGND sg13g2_fill_1
XFILLER_40_618 VPWR VGND sg13g2_decap_8
XFILLER_40_607 VPWR VGND sg13g2_fill_2
XFILLER_36_1001 VPWR VGND sg13g2_decap_8
X_5985_ net30 VGND VPWR _0035_ s0.shift_out\[19\][0] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_40_629 VPWR VGND sg13g2_fill_2
X_4936_ _0649_ _0650_ _0073_ VPWR VGND sg13g2_nor2_1
X_4867_ VGND VPWR _0500_ _0584_ _0585_ net1149 sg13g2_a21oi_1
XFILLER_21_843 VPWR VGND sg13g2_decap_8
X_3818_ net950 net1057 _2207_ VPWR VGND sg13g2_nor2b_1
X_4798_ net1148 VPWR _0525_ VGND net1228 net1137 sg13g2_o21ai_1
X_3749_ VGND VPWR _2146_ _2139_ net1234 sg13g2_or2_1
XFILLER_21_58 VPWR VGND sg13g2_fill_1
X_5419_ s0.data_out\[12\]\[6\] s0.data_out\[11\]\[6\] net1098 _1088_ VPWR VGND sg13g2_mux2_1
XFILLER_0_747 VPWR VGND sg13g2_decap_8
XFILLER_46_44 VPWR VGND sg13g2_decap_8
XFILLER_44_913 VPWR VGND sg13g2_decap_8
XFILLER_28_453 VPWR VGND sg13g2_fill_1
XFILLER_16_659 VPWR VGND sg13g2_decap_4
XFILLER_28_486 VPWR VGND sg13g2_fill_2
XFILLER_43_478 VPWR VGND sg13g2_decap_8
XFILLER_7_27 VPWR VGND sg13g2_fill_2
XFILLER_7_379 VPWR VGND sg13g2_decap_4
Xfanout1320 net1322 net1320 VPWR VGND sg13g2_buf_8
Xfanout1331 net1349 net1331 VPWR VGND sg13g2_buf_2
Xfanout1342 net1348 net1342 VPWR VGND sg13g2_buf_8
XFILLER_47_773 VPWR VGND sg13g2_decap_8
XFILLER_35_957 VPWR VGND sg13g2_decap_8
XFILLER_19_497 VPWR VGND sg13g2_fill_1
X_5770_ _1398_ VPWR _1399_ VGND net1343 net385 sg13g2_o21ai_1
XFILLER_22_629 VPWR VGND sg13g2_decap_8
X_4721_ _0450_ _0453_ net1306 _0454_ VPWR VGND sg13g2_nand3_1
XFILLER_21_139 VPWR VGND sg13g2_decap_8
X_4652_ _0393_ net1165 net582 VPWR VGND sg13g2_nand2_1
X_3603_ VPWR VGND _1945_ net1284 _2010_ net1275 _2012_ _2007_ sg13g2_a221oi_1
X_4583_ net1169 VPWR _0329_ VGND _0327_ _0328_ sg13g2_o21ai_1
X_3534_ VPWR _0214_ _1950_ VGND sg13g2_inv_1
XFILLER_6_390 VPWR VGND sg13g2_decap_8
X_3465_ VGND VPWR net990 _1885_ _1886_ _1842_ sg13g2_a21oi_1
X_5204_ _0889_ _0892_ net1332 _0893_ VPWR VGND sg13g2_nand3_1
X_3396_ _1825_ _1826_ _0200_ VPWR VGND sg13g2_nor2_1
X_6184_ net87 VGND VPWR _0234_ s0.shift_out\[3\][0] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_5135_ _0827_ net1112 _0787_ _0828_ VPWR VGND sg13g2_a21o_1
X_5066_ _0767_ _0768_ _0769_ VPWR VGND sg13g2_nor2b_1
X_4017_ net1247 _2387_ _2390_ VPWR VGND sg13g2_nor2_1
XFILLER_41_905 VPWR VGND sg13g2_decap_8
X_5968_ net48 VGND VPWR _0018_ s0.data_out\[20\]\[3\] clknet_leaf_36_clk sg13g2_dfrbpq_2
X_4919_ _0626_ VPWR _0636_ VGND _0625_ _0631_ sg13g2_o21ai_1
XFILLER_21_640 VPWR VGND sg13g2_decap_8
X_5899_ net1342 VPWR _1516_ VGND net918 _1515_ sg13g2_o21ai_1
XFILLER_20_161 VPWR VGND sg13g2_decap_4
XFILLER_32_79 VPWR VGND sg13g2_decap_8
XFILLER_5_839 VPWR VGND sg13g2_decap_8
XFILLER_0_544 VPWR VGND sg13g2_decap_8
XFILLER_28_272 VPWR VGND sg13g2_decap_8
XFILLER_16_434 VPWR VGND sg13g2_fill_2
XFILLER_32_905 VPWR VGND sg13g2_fill_2
XFILLER_7_154 VPWR VGND sg13g2_fill_1
XFILLER_4_872 VPWR VGND sg13g2_decap_8
X_3250_ _1695_ _1691_ _1692_ _1694_ VPWR VGND sg13g2_and3_1
XFILLER_26_1022 VPWR VGND sg13g2_decap_8
X_3181_ _1629_ net539 net1020 VPWR VGND sg13g2_nand2b_1
Xfanout1150 net338 net1150 VPWR VGND sg13g2_buf_2
XFILLER_21_4 VPWR VGND sg13g2_decap_8
XFILLER_39_548 VPWR VGND sg13g2_fill_2
Xfanout1161 net1162 net1161 VPWR VGND sg13g2_buf_8
Xfanout1183 net1185 net1183 VPWR VGND sg13g2_buf_8
Xfanout1172 net1173 net1172 VPWR VGND sg13g2_buf_8
Xfanout1194 net333 net1194 VPWR VGND sg13g2_buf_2
X_5822_ _1448_ _1444_ _1447_ VPWR VGND sg13g2_nand2_1
XFILLER_22_404 VPWR VGND sg13g2_decap_8
XFILLER_22_459 VPWR VGND sg13g2_decap_4
X_5753_ _1380_ _1383_ net1341 _1384_ VPWR VGND sg13g2_nand3_1
XFILLER_34_297 VPWR VGND sg13g2_fill_2
X_6221__71 VPWR VGND net71 sg13g2_tiehi
X_4704_ net1304 VPWR _0439_ VGND net924 _0438_ sg13g2_o21ai_1
XFILLER_31_971 VPWR VGND sg13g2_decap_8
XFILLER_33_1004 VPWR VGND sg13g2_decap_8
XFILLER_30_481 VPWR VGND sg13g2_decap_8
X_5684_ VGND VPWR net1040 _1328_ _1329_ _1270_ sg13g2_a21oi_1
X_4635_ VGND VPWR net1155 _0375_ _0376_ _0328_ sg13g2_a21oi_1
X_4566_ VGND VPWR net1156 s0.data_out\[17\]\[1\] _0314_ _0313_ sg13g2_a21oi_1
X_3517_ _1936_ _1935_ _1934_ VPWR VGND sg13g2_nand2b_1
X_4497_ VGND VPWR _2756_ _2811_ _2813_ net1275 sg13g2_a21oi_1
X_3448_ net985 net1050 _1871_ VPWR VGND sg13g2_nor2b_1
X_5995__291 VPWR VGND net291 sg13g2_tiehi
X_6167_ net105 VGND VPWR _0217_ s0.data_out\[4\]\[3\] clknet_leaf_14_clk sg13g2_dfrbpq_2
X_3379_ _1802_ VPWR _1812_ VGND _1808_ _1809_ sg13g2_o21ai_1
XFILLER_40_1008 VPWR VGND sg13g2_decap_8
X_5118_ _0813_ net597 net1132 VPWR VGND sg13g2_nand2b_1
X_6098_ net180 VGND VPWR _0148_ s0.data_new_delayed\[4\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_38_592 VPWR VGND sg13g2_fill_1
X_5049_ _0754_ net1215 _0745_ VPWR VGND sg13g2_xnor2_1
XFILLER_13_426 VPWR VGND sg13g2_fill_2
XFILLER_25_297 VPWR VGND sg13g2_decap_4
XFILLER_22_971 VPWR VGND sg13g2_decap_8
XFILLER_4_39 VPWR VGND sg13g2_fill_1
XFILLER_0_352 VPWR VGND sg13g2_fill_1
XFILLER_1_886 VPWR VGND sg13g2_decap_8
XFILLER_49_835 VPWR VGND sg13g2_decap_8
XFILLER_48_378 VPWR VGND sg13g2_decap_4
XFILLER_44_540 VPWR VGND sg13g2_fill_2
XFILLER_17_743 VPWR VGND sg13g2_decap_8
XFILLER_31_278 VPWR VGND sg13g2_fill_1
XFILLER_9_964 VPWR VGND sg13g2_decap_8
X_4420_ _2746_ _2743_ _2745_ VPWR VGND sg13g2_nand2_1
X_4351_ _2680_ VPWR _2681_ VGND _2676_ _2679_ sg13g2_o21ai_1
X_4282_ VGND VPWR _2622_ net1208 net306 sg13g2_or2_1
X_3302_ VPWR _0193_ _1739_ VGND sg13g2_inv_1
X_3233_ net1250 _1676_ _1678_ VPWR VGND sg13g2_nor2_1
X_6021_ net263 VGND VPWR _0071_ s0.shift_out\[16\][0] clknet_leaf_32_clk sg13g2_dfrbpq_1
XFILLER_39_312 VPWR VGND sg13g2_fill_2
X_3164_ VPWR _0180_ _1614_ VGND sg13g2_inv_1
XFILLER_27_529 VPWR VGND sg13g2_decap_8
XFILLER_23_702 VPWR VGND sg13g2_fill_1
XFILLER_35_595 VPWR VGND sg13g2_decap_8
X_3997_ _2369_ net943 _2342_ _2370_ VPWR VGND sg13g2_a21o_1
X_5805_ _1431_ net1035 _1430_ VPWR VGND sg13g2_nand2b_1
X_5736_ net1035 VPWR _1369_ VGND _1367_ _1368_ sg13g2_o21ai_1
XFILLER_31_790 VPWR VGND sg13g2_fill_2
X_5667_ _1312_ _1311_ net1265 _1297_ net1270 VPWR VGND sg13g2_a22oi_1
X_4618_ VPWR _0046_ net580 VGND sg13g2_inv_1
X_5598_ net1077 VPWR _1250_ VGND _1248_ _1249_ sg13g2_o21ai_1
X_4549_ net925 VPWR _0300_ VGND net375 net1177 sg13g2_o21ai_1
Xfanout932 _2455_ net932 VPWR VGND sg13g2_buf_8
Xfanout943 net944 net943 VPWR VGND sg13g2_buf_8
X_6219_ net97 VGND VPWR _0269_ s0.data_out\[0\]\[7\] clknet_leaf_9_clk sg13g2_dfrbpq_2
Xfanout921 _2464_ net921 VPWR VGND sg13g2_buf_8
Xfanout954 s0.shift_out\[1\][0] net954 VPWR VGND sg13g2_buf_8
Xfanout976 net979 net976 VPWR VGND sg13g2_buf_8
Xfanout965 net968 net965 VPWR VGND sg13g2_buf_8
Xfanout998 net999 net998 VPWR VGND sg13g2_buf_8
Xfanout987 net989 net987 VPWR VGND sg13g2_buf_8
XFILLER_46_838 VPWR VGND sg13g2_decap_8
XFILLER_45_359 VPWR VGND sg13g2_decap_8
XFILLER_41_510 VPWR VGND sg13g2_decap_4
XFILLER_16_1021 VPWR VGND sg13g2_decap_8
XFILLER_6_912 VPWR VGND sg13g2_decap_8
XFILLER_10_996 VPWR VGND sg13g2_decap_8
XFILLER_6_989 VPWR VGND sg13g2_decap_8
XFILLER_5_433 VPWR VGND sg13g2_fill_2
XFILLER_5_488 VPWR VGND sg13g2_fill_2
XFILLER_49_632 VPWR VGND sg13g2_decap_8
XFILLER_1_683 VPWR VGND sg13g2_decap_8
XFILLER_37_849 VPWR VGND sg13g2_decap_8
Xheichips25_top_sorter_295 VPWR VGND uio_oe[2] sg13g2_tiehi
X_3920_ net942 s0.data_out\[0\]\[1\] _2300_ VPWR VGND sg13g2_and2_1
XFILLER_45_893 VPWR VGND sg13g2_decap_8
XFILLER_32_510 VPWR VGND sg13g2_fill_1
XFILLER_20_716 VPWR VGND sg13g2_decap_8
X_3851_ s0.data_out\[2\]\[1\] s0.data_out\[1\]\[1\] net955 _2236_ VPWR VGND sg13g2_mux2_1
X_3782_ net1218 _2170_ _0237_ VPWR VGND sg13g2_nor2_1
XFILLER_20_727 VPWR VGND sg13g2_fill_1
XFILLER_9_750 VPWR VGND sg13g2_decap_8
X_5521_ VGND VPWR _1179_ net540 net1345 sg13g2_or2_1
X_5452_ VGND VPWR _1119_ _1118_ _1117_ sg13g2_or2_1
X_4403_ _2729_ _2730_ _2731_ VPWR VGND sg13g2_nor2_1
X_5383_ _1053_ VPWR _1054_ VGND _1049_ _1052_ sg13g2_o21ai_1
X_4334_ _2662_ _2665_ net1289 _2666_ VPWR VGND sg13g2_nand3_1
X_6004_ net281 VGND VPWR _0054_ s0.data_out\[17\]\[3\] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_4265_ VGND VPWR net1204 _2604_ _2605_ _2547_ sg13g2_a21oi_1
XFILLER_39_131 VPWR VGND sg13g2_fill_2
X_4196_ net1216 _2540_ _2541_ VPWR VGND sg13g2_nor2_1
X_5992__294 VPWR VGND net294 sg13g2_tiehi
X_3216_ _1595_ VPWR _1661_ VGND net917 _1660_ sg13g2_o21ai_1
X_3147_ _1599_ VPWR _1600_ VGND net1327 net391 sg13g2_o21ai_1
XFILLER_42_318 VPWR VGND sg13g2_decap_4
XFILLER_39_1021 VPWR VGND sg13g2_decap_8
XFILLER_23_565 VPWR VGND sg13g2_fill_2
X_6179__92 VPWR VGND net92 sg13g2_tiehi
XFILLER_40_35 VPWR VGND sg13g2_decap_4
X_5719_ _1354_ VPWR _1355_ VGND net1028 _1348_ sg13g2_o21ai_1
XFILLER_3_915 VPWR VGND sg13g2_decap_8
XFILLER_2_414 VPWR VGND sg13g2_fill_2
Xhold271 s0.data_out\[19\]\[3\] VPWR VGND net567 sg13g2_dlygate4sd3_1
XFILLER_2_425 VPWR VGND sg13g2_fill_2
Xhold260 s0.data_out\[12\]\[4\] VPWR VGND net556 sg13g2_dlygate4sd3_1
Xhold293 s0.data_out\[7\]\[5\] VPWR VGND net589 sg13g2_dlygate4sd3_1
Xhold282 _0826_ VPWR VGND net578 sg13g2_dlygate4sd3_1
XFILLER_45_112 VPWR VGND sg13g2_fill_2
XFILLER_14_510 VPWR VGND sg13g2_fill_1
XFILLER_14_554 VPWR VGND sg13g2_fill_1
XFILLER_14_565 VPWR VGND sg13g2_decap_8
XFILLER_14_598 VPWR VGND sg13g2_fill_2
XFILLER_5_241 VPWR VGND sg13g2_fill_1
X_4050_ net1218 _2414_ _2415_ VPWR VGND sg13g2_nor2_1
XFILLER_37_657 VPWR VGND sg13g2_fill_2
XFILLER_37_635 VPWR VGND sg13g2_fill_1
XFILLER_25_808 VPWR VGND sg13g2_decap_4
XFILLER_37_679 VPWR VGND sg13g2_fill_1
XFILLER_45_690 VPWR VGND sg13g2_decap_8
X_4952_ _0663_ VPWR _0664_ VGND net1318 net431 sg13g2_o21ai_1
XFILLER_18_893 VPWR VGND sg13g2_fill_1
X_3903_ _2284_ VPWR _2286_ VGND s0.was_valid_out\[0\][0] net947 sg13g2_o21ai_1
X_4883_ VGND VPWR net1134 _0599_ _0600_ _0538_ sg13g2_a21oi_1
XFILLER_17_392 VPWR VGND sg13g2_decap_8
XFILLER_33_863 VPWR VGND sg13g2_decap_4
X_3834_ VGND VPWR net953 s0.data_out\[1\]\[6\] _2221_ _2220_ sg13g2_a21oi_1
XFILLER_20_502 VPWR VGND sg13g2_fill_1
X_3765_ _2147_ _2155_ _2156_ _2162_ VPWR VGND sg13g2_nor3_1
X_3696_ _2096_ net349 net977 VPWR VGND sg13g2_nand2b_1
X_5504_ net1345 VPWR _1164_ VGND net939 _1163_ sg13g2_o21ai_1
X_6176__95 VPWR VGND net95 sg13g2_tiehi
X_5435_ _1104_ net1251 _1103_ VPWR VGND sg13g2_nand2_1
XFILLER_0_929 VPWR VGND sg13g2_decap_8
X_5366_ VGND VPWR _1039_ net556 net1337 sg13g2_or2_1
X_4317_ net1286 VPWR _2651_ VGND net931 _2650_ sg13g2_o21ai_1
X_5297_ _0978_ net1109 s0.data_out\[12\]\[4\] VPWR VGND sg13g2_nand2_1
X_4248_ _2588_ net1260 _2587_ VPWR VGND sg13g2_nand2_1
XFILLER_19_36 VPWR VGND sg13g2_decap_8
X_4179_ _2523_ _2525_ net1285 _2526_ VPWR VGND sg13g2_nand3_1
XFILLER_16_808 VPWR VGND sg13g2_decap_4
XFILLER_27_112 VPWR VGND sg13g2_fill_2
XFILLER_15_329 VPWR VGND sg13g2_fill_1
Xclkbuf_3_3__f_clk clknet_0_clk clknet_3_3__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_11_546 VPWR VGND sg13g2_decap_8
XFILLER_7_517 VPWR VGND sg13g2_decap_8
XFILLER_3_712 VPWR VGND sg13g2_decap_8
XFILLER_2_200 VPWR VGND sg13g2_decap_8
XFILLER_3_789 VPWR VGND sg13g2_decap_8
XFILLER_2_299 VPWR VGND sg13g2_fill_2
XFILLER_47_955 VPWR VGND sg13g2_decap_8
XFILLER_18_167 VPWR VGND sg13g2_decap_4
XFILLER_34_605 VPWR VGND sg13g2_decap_8
XFILLER_18_178 VPWR VGND sg13g2_decap_4
XFILLER_42_693 VPWR VGND sg13g2_decap_4
XFILLER_41_181 VPWR VGND sg13g2_fill_2
XFILLER_30_855 VPWR VGND sg13g2_decap_4
X_3550_ VPWR _0216_ net534 VGND sg13g2_inv_1
X_5220_ _0903_ _0906_ net1332 _0907_ VPWR VGND sg13g2_nand3_1
X_3481_ _1901_ VPWR _1902_ VGND _1895_ _1896_ sg13g2_o21ai_1
X_5151_ _0793_ _0843_ _0844_ VPWR VGND sg13g2_and2_1
X_5082_ net1333 VPWR _0782_ VGND net937 _0781_ sg13g2_o21ai_1
X_4102_ _2461_ net1171 VPWR VGND sg13g2_inv_2
XFILLER_38_933 VPWR VGND sg13g2_decap_8
X_4033_ net377 net1218 _2401_ _0262_ VPWR VGND sg13g2_a21o_1
XFILLER_49_270 VPWR VGND sg13g2_fill_1
XFILLER_25_627 VPWR VGND sg13g2_fill_2
X_5984_ net31 VGND VPWR _0034_ s0.data_out\[19\]\[7\] clknet_leaf_0_clk sg13g2_dfrbpq_2
X_4935_ net1319 VPWR _0650_ VGND net381 _0645_ sg13g2_o21ai_1
X_4866_ _0584_ net554 net1152 VPWR VGND sg13g2_nand2b_1
XFILLER_21_866 VPWR VGND sg13g2_fill_2
XFILLER_32_192 VPWR VGND sg13g2_fill_2
X_3817_ net950 s0.data_out\[1\]\[4\] _2206_ VPWR VGND sg13g2_and2_1
X_4797_ net1319 net310 _0060_ VPWR VGND sg13g2_and2_1
XFILLER_21_888 VPWR VGND sg13g2_fill_1
X_3748_ net1241 _2143_ _2145_ VPWR VGND sg13g2_nor2_1
XFILLER_20_387 VPWR VGND sg13g2_fill_1
X_3679_ VPWR _0228_ _2081_ VGND sg13g2_inv_1
X_5418_ _1087_ net1097 net527 VPWR VGND sg13g2_nand2_1
XFILLER_0_726 VPWR VGND sg13g2_decap_8
X_5349_ net1334 VPWR _1024_ VGND net938 _1023_ sg13g2_o21ai_1
XFILLER_43_1028 VPWR VGND sg13g2_fill_1
XFILLER_43_1017 VPWR VGND sg13g2_decap_8
XFILLER_16_605 VPWR VGND sg13g2_fill_2
XFILLER_29_988 VPWR VGND sg13g2_decap_8
XFILLER_44_969 VPWR VGND sg13g2_decap_8
XFILLER_30_118 VPWR VGND sg13g2_decap_8
XFILLER_31_619 VPWR VGND sg13g2_fill_2
X_6027__256 VPWR VGND net256 sg13g2_tiehi
XFILLER_7_314 VPWR VGND sg13g2_fill_1
XFILLER_7_303 VPWR VGND sg13g2_fill_1
XFILLER_12_877 VPWR VGND sg13g2_decap_8
XFILLER_8_848 VPWR VGND sg13g2_fill_2
XFILLER_3_564 VPWR VGND sg13g2_decap_4
XFILLER_30_9 VPWR VGND sg13g2_fill_1
Xfanout1332 net1333 net1332 VPWR VGND sg13g2_buf_8
Xfanout1321 net1322 net1321 VPWR VGND sg13g2_buf_2
Xfanout1310 net1316 net1310 VPWR VGND sg13g2_buf_8
Xfanout1343 net1348 net1343 VPWR VGND sg13g2_buf_1
X_6034__249 VPWR VGND net249 sg13g2_tiehi
XFILLER_47_752 VPWR VGND sg13g2_decap_8
XFILLER_46_251 VPWR VGND sg13g2_fill_1
XFILLER_46_295 VPWR VGND sg13g2_fill_1
XFILLER_21_118 VPWR VGND sg13g2_decap_4
X_4720_ net1161 VPWR _0453_ VGND _0451_ _0452_ sg13g2_o21ai_1
X_4651_ _0391_ _0389_ _0392_ VPWR VGND _0390_ sg13g2_nand3b_1
X_3602_ _2003_ VPWR _2011_ VGND net1275 _2007_ sg13g2_o21ai_1
X_4582_ net1156 net1061 _0328_ VPWR VGND sg13g2_nor2b_1
X_3533_ _1949_ VPWR _1950_ VGND net1308 net440 sg13g2_o21ai_1
XFILLER_42_0 VPWR VGND sg13g2_decap_8
X_3464_ _1884_ net981 _1843_ _1885_ VPWR VGND sg13g2_a21o_1
X_6183_ net88 VGND VPWR _0233_ s0.data_out\[3\]\[7\] clknet_leaf_12_clk sg13g2_dfrbpq_2
X_5203_ net1116 VPWR _0892_ VGND _0890_ _0891_ sg13g2_o21ai_1
X_3395_ net1313 VPWR _1826_ VGND net383 _1821_ sg13g2_o21ai_1
X_5134_ s0.data_out\[14\]\[2\] s0.data_out\[13\]\[2\] net1119 _0827_ VPWR VGND sg13g2_mux2_1
XFILLER_29_218 VPWR VGND sg13g2_fill_2
X_5065_ net937 VPWR _0768_ VGND net346 net1132 sg13g2_o21ai_1
X_4016_ VGND VPWR _2389_ _2365_ net1261 sg13g2_or2_1
X_5967_ net49 VGND VPWR _0017_ s0.data_out\[20\]\[2\] clknet_leaf_0_clk sg13g2_dfrbpq_2
XFILLER_12_118 VPWR VGND sg13g2_fill_1
X_4918_ _0634_ VPWR _0635_ VGND _0603_ _0609_ sg13g2_o21ai_1
Xclkbuf_leaf_32_clk clknet_3_4__leaf_clk clknet_leaf_32_clk VPWR VGND sg13g2_buf_8
XFILLER_33_490 VPWR VGND sg13g2_decap_4
XFILLER_34_991 VPWR VGND sg13g2_decap_8
X_5898_ VGND VPWR net1016 s0.data_out\[7\]\[5\] _1515_ _1514_ sg13g2_a21oi_1
X_4849_ VPWR _0067_ _0569_ VGND sg13g2_inv_1
XFILLER_21_685 VPWR VGND sg13g2_decap_4
XFILLER_32_69 VPWR VGND sg13g2_fill_1
XFILLER_5_818 VPWR VGND sg13g2_decap_8
XFILLER_0_523 VPWR VGND sg13g2_decap_8
XFILLER_48_527 VPWR VGND sg13g2_decap_8
XFILLER_29_763 VPWR VGND sg13g2_fill_1
XFILLER_44_722 VPWR VGND sg13g2_fill_2
XFILLER_28_295 VPWR VGND sg13g2_fill_2
XFILLER_44_788 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_23_clk clknet_3_4__leaf_clk clknet_leaf_23_clk VPWR VGND sg13g2_buf_8
XFILLER_8_612 VPWR VGND sg13g2_decap_8
XFILLER_40_994 VPWR VGND sg13g2_decap_8
X_6040__242 VPWR VGND net242 sg13g2_tiehi
XFILLER_4_851 VPWR VGND sg13g2_decap_8
XFILLER_26_1001 VPWR VGND sg13g2_decap_8
X_3180_ VPWR _0182_ _1628_ VGND sg13g2_inv_1
Xfanout1140 net336 net1140 VPWR VGND sg13g2_buf_8
XFILLER_39_538 VPWR VGND sg13g2_fill_1
Xfanout1162 s0.shift_out\[17\][0] net1162 VPWR VGND sg13g2_buf_8
Xfanout1151 net1154 net1151 VPWR VGND sg13g2_buf_8
XFILLER_14_4 VPWR VGND sg13g2_fill_2
Xfanout1173 s0.shift_out\[18\][0] net1173 VPWR VGND sg13g2_buf_8
Xfanout1184 net1185 net1184 VPWR VGND sg13g2_buf_1
Xfanout1195 net1196 net1195 VPWR VGND sg13g2_buf_8
XFILLER_47_571 VPWR VGND sg13g2_decap_8
XFILLER_35_700 VPWR VGND sg13g2_fill_2
XFILLER_35_744 VPWR VGND sg13g2_decap_8
X_5821_ VGND VPWR _1447_ _1439_ net1237 sg13g2_or2_1
XFILLER_22_427 VPWR VGND sg13g2_fill_2
XFILLER_22_438 VPWR VGND sg13g2_fill_1
X_5752_ net1035 VPWR _1383_ VGND _1381_ _1382_ sg13g2_o21ai_1
Xclkbuf_leaf_14_clk clknet_3_3__leaf_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
X_4703_ VGND VPWR net1144 net422 _0438_ _0437_ sg13g2_a21oi_1
XFILLER_31_950 VPWR VGND sg13g2_decap_8
X_5683_ s0.data_out\[10\]\[4\] s0.data_out\[9\]\[4\] net1043 _1328_ VPWR VGND sg13g2_mux2_1
X_4634_ s0.data_out\[18\]\[3\] s0.data_out\[17\]\[3\] net1163 _0375_ VPWR VGND sg13g2_mux2_1
X_4565_ net1155 net1072 _0313_ VPWR VGND sg13g2_nor2b_1
X_3516_ _1935_ net1222 net977 VPWR VGND sg13g2_nand2_1
X_4496_ _2756_ _2811_ net1275 _2812_ VPWR VGND sg13g2_nand3_1
X_3447_ VGND VPWR _1791_ _1869_ _1870_ net994 sg13g2_a21oi_1
X_6166_ net106 VGND VPWR _0216_ s0.data_out\[4\]\[2\] clknet_leaf_5_clk sg13g2_dfrbpq_2
X_3378_ _1807_ _1808_ _1786_ _1811_ VPWR VGND _1810_ sg13g2_nand4_1
X_5117_ VPWR _0092_ net549 VGND sg13g2_inv_1
X_6097_ net181 VGND VPWR _0147_ s0.data_new_delayed\[3\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_5048_ VGND VPWR _0687_ _0750_ _0753_ net1250 sg13g2_a21oi_1
XFILLER_38_582 VPWR VGND sg13g2_fill_1
XFILLER_26_700 VPWR VGND sg13g2_decap_8
XFILLER_41_725 VPWR VGND sg13g2_decap_8
XFILLER_25_254 VPWR VGND sg13g2_fill_1
XFILLER_22_950 VPWR VGND sg13g2_decap_8
X_6024__259 VPWR VGND net259 sg13g2_tiehi
XFILLER_4_29 VPWR VGND sg13g2_fill_1
XFILLER_49_814 VPWR VGND sg13g2_decap_8
XFILLER_1_865 VPWR VGND sg13g2_decap_8
XFILLER_0_386 VPWR VGND sg13g2_decap_8
XFILLER_31_213 VPWR VGND sg13g2_fill_1
XFILLER_9_943 VPWR VGND sg13g2_decap_8
XFILLER_8_486 VPWR VGND sg13g2_fill_1
X_4350_ VGND VPWR _2680_ net592 net1288 sg13g2_or2_1
X_3301_ _1738_ VPWR _1739_ VGND net1324 net454 sg13g2_o21ai_1
X_4281_ _2621_ net1223 net1292 VPWR VGND sg13g2_nand2_1
X_3232_ _1677_ _1676_ net1250 _1672_ net1258 VPWR VGND sg13g2_a22oi_1
X_6020_ net264 VGND VPWR _0070_ s0.data_out\[16\]\[7\] clknet_leaf_34_clk sg13g2_dfrbpq_2
Xclkbuf_leaf_3_clk clknet_3_1__leaf_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
X_3163_ _1613_ VPWR _1614_ VGND net1324 net467 sg13g2_o21ai_1
XFILLER_39_357 VPWR VGND sg13g2_fill_1
XFILLER_35_563 VPWR VGND sg13g2_fill_1
XFILLER_22_202 VPWR VGND sg13g2_fill_1
X_5804_ VGND VPWR net1030 _1429_ _1430_ _1382_ sg13g2_a21oi_1
X_3996_ s0.data_out\[1\]\[7\] s0.data_out\[0\]\[7\] net948 _2369_ VPWR VGND sg13g2_mux2_1
X_5735_ net1030 net1071 _1368_ VPWR VGND sg13g2_nor2b_1
X_5666_ _1261_ _1310_ _1311_ VPWR VGND sg13g2_and2_1
X_4617_ _0358_ VPWR _0359_ VGND _0354_ _0357_ sg13g2_o21ai_1
X_5597_ net1036 net1071 _1249_ VPWR VGND sg13g2_nor2b_1
XFILLER_2_629 VPWR VGND sg13g2_decap_8
X_4548_ VGND VPWR _0299_ net1166 net375 sg13g2_or2_1
XFILLER_8_9 VPWR VGND sg13g2_decap_8
X_4479_ VPWR _0033_ net552 VGND sg13g2_inv_1
Xfanout933 _2455_ net933 VPWR VGND sg13g2_buf_1
X_6218_ net110 VGND VPWR _0268_ s0.data_out\[0\]\[6\] clknet_leaf_8_clk sg13g2_dfrbpq_2
Xfanout922 _2463_ net922 VPWR VGND sg13g2_buf_8
Xfanout977 net979 net977 VPWR VGND sg13g2_buf_8
Xfanout944 net945 net944 VPWR VGND sg13g2_buf_8
Xfanout966 net968 net966 VPWR VGND sg13g2_buf_8
XFILLER_38_13 VPWR VGND sg13g2_decap_8
Xfanout955 net958 net955 VPWR VGND sg13g2_buf_8
X_6149_ net125 VGND VPWR _0199_ s0.genblk1\[5\].modules.bubble clknet_leaf_12_clk
+ sg13g2_dfrbpq_1
XFILLER_46_817 VPWR VGND sg13g2_decap_8
Xfanout988 net989 net988 VPWR VGND sg13g2_buf_8
Xfanout999 s0.valid_out\[5\][0] net999 VPWR VGND sg13g2_buf_8
XFILLER_18_519 VPWR VGND sg13g2_decap_8
XFILLER_38_390 VPWR VGND sg13g2_fill_1
XFILLER_26_530 VPWR VGND sg13g2_decap_4
XFILLER_14_758 VPWR VGND sg13g2_decap_8
XFILLER_14_769 VPWR VGND sg13g2_fill_2
XFILLER_16_1000 VPWR VGND sg13g2_decap_8
XFILLER_41_599 VPWR VGND sg13g2_decap_4
XFILLER_41_577 VPWR VGND sg13g2_fill_2
XFILLER_9_239 VPWR VGND sg13g2_decap_4
XFILLER_5_412 VPWR VGND sg13g2_fill_2
XFILLER_10_975 VPWR VGND sg13g2_decap_8
XFILLER_6_968 VPWR VGND sg13g2_decap_8
XFILLER_5_445 VPWR VGND sg13g2_fill_2
XFILLER_1_662 VPWR VGND sg13g2_decap_8
XFILLER_49_611 VPWR VGND sg13g2_decap_8
XFILLER_0_172 VPWR VGND sg13g2_fill_2
XFILLER_48_132 VPWR VGND sg13g2_fill_1
XFILLER_49_688 VPWR VGND sg13g2_decap_8
XFILLER_37_839 VPWR VGND sg13g2_decap_4
XFILLER_36_338 VPWR VGND sg13g2_decap_8
Xheichips25_top_sorter_296 VPWR VGND uio_oe[5] sg13g2_tiehi
XFILLER_45_872 VPWR VGND sg13g2_decap_8
X_3850_ VGND VPWR _2235_ _2234_ net1268 sg13g2_or2_1
X_3781_ VGND VPWR _2171_ _2174_ _0236_ _2175_ sg13g2_a21oi_1
XFILLER_13_780 VPWR VGND sg13g2_fill_1
X_6188__82 VPWR VGND net82 sg13g2_tiehi
X_5520_ net1344 VPWR _1178_ VGND _2448_ _1177_ sg13g2_o21ai_1
XFILLER_9_773 VPWR VGND sg13g2_decap_8
XFILLER_9_784 VPWR VGND sg13g2_fill_1
X_5451_ net1094 _0997_ _1118_ VPWR VGND sg13g2_nor2_1
X_4402_ net1260 _2706_ _2730_ VPWR VGND sg13g2_nor2_1
X_5382_ VGND VPWR _1053_ net588 net1336 sg13g2_or2_1
X_4333_ net1196 VPWR _2665_ VGND _2663_ _2664_ sg13g2_o21ai_1
X_4264_ _2603_ net1195 _2543_ _2604_ VPWR VGND sg13g2_a21o_1
X_6003_ net282 VGND VPWR _0053_ s0.data_out\[17\]\[2\] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_3215_ VGND VPWR net1001 _1659_ _1660_ _1597_ sg13g2_a21oi_1
X_4195_ net1202 _2538_ _2539_ _2540_ VPWR VGND sg13g2_nor3_1
XFILLER_28_806 VPWR VGND sg13g2_fill_1
X_3146_ _1595_ _1598_ net1327 _1599_ VPWR VGND sg13g2_nand3_1
XFILLER_27_316 VPWR VGND sg13g2_fill_1
XFILLER_39_1000 VPWR VGND sg13g2_decap_8
XFILLER_35_360 VPWR VGND sg13g2_decap_8
XFILLER_35_393 VPWR VGND sg13g2_decap_4
XFILLER_11_706 VPWR VGND sg13g2_decap_8
XFILLER_23_577 VPWR VGND sg13g2_decap_4
X_5718_ net920 VPWR _1354_ VGND net398 net1042 sg13g2_o21ai_1
X_3979_ VGND VPWR net942 _2351_ _2352_ _2301_ sg13g2_a21oi_1
X_5649_ VPWR _0142_ net532 VGND sg13g2_inv_1
Xhold261 s0.data_out\[6\]\[6\] VPWR VGND net557 sg13g2_dlygate4sd3_1
XFILLER_6_6 VPWR VGND sg13g2_fill_1
Xhold250 s0.data_out\[16\]\[6\] VPWR VGND net546 sg13g2_dlygate4sd3_1
Xhold294 s0.data_out\[1\]\[6\] VPWR VGND net590 sg13g2_dlygate4sd3_1
Xhold283 s0.data_out\[18\]\[7\] VPWR VGND net579 sg13g2_dlygate4sd3_1
Xhold272 s0.data_out\[11\]\[2\] VPWR VGND net568 sg13g2_dlygate4sd3_1
X_6169__103 VPWR VGND net103 sg13g2_tiehi
XFILLER_45_124 VPWR VGND sg13g2_fill_1
XFILLER_34_809 VPWR VGND sg13g2_fill_1
XFILLER_45_168 VPWR VGND sg13g2_fill_1
XFILLER_14_522 VPWR VGND sg13g2_fill_2
XFILLER_27_894 VPWR VGND sg13g2_fill_1
XFILLER_41_374 VPWR VGND sg13g2_fill_2
XFILLER_41_352 VPWR VGND sg13g2_decap_4
XFILLER_6_776 VPWR VGND sg13g2_decap_8
XFILLER_5_297 VPWR VGND sg13g2_fill_1
XFILLER_7_1020 VPWR VGND sg13g2_decap_8
XFILLER_49_485 VPWR VGND sg13g2_decap_8
XFILLER_18_861 VPWR VGND sg13g2_fill_1
X_4951_ _0659_ _0662_ net1318 _0663_ VPWR VGND sg13g2_nand3_1
X_3902_ VGND VPWR net928 _2167_ _2285_ _2284_ sg13g2_a21oi_1
X_4882_ s0.data_out\[16\]\[0\] s0.data_out\[15\]\[0\] net1141 _0599_ VPWR VGND sg13g2_mux2_1
X_3833_ net953 net1049 _2220_ VPWR VGND sg13g2_nor2b_1
XFILLER_32_385 VPWR VGND sg13g2_fill_1
X_3764_ _2147_ _2159_ _2160_ _2161_ VPWR VGND sg13g2_or3_1
X_5503_ VGND VPWR net1080 net481 _1163_ _1162_ sg13g2_a21oi_1
X_3695_ VPWR _0230_ _2095_ VGND sg13g2_inv_1
X_5434_ VGND VPWR net1105 _1102_ _1103_ _1042_ sg13g2_a21oi_1
XFILLER_0_908 VPWR VGND sg13g2_decap_8
X_5365_ net1337 VPWR _1038_ VGND net938 _1037_ sg13g2_o21ai_1
X_4316_ VGND VPWR net1179 net475 _2650_ _2649_ sg13g2_a21oi_1
X_5296_ _0977_ _0973_ _0974_ _0976_ VPWR VGND sg13g2_and3_1
X_4247_ VGND VPWR net1203 _2586_ _2587_ _2540_ sg13g2_a21oi_1
X_4178_ _2524_ VPWR _2525_ VGND net1206 s0.data_out\[20\]\[1\] sg13g2_o21ai_1
XFILLER_28_625 VPWR VGND sg13g2_fill_2
X_3129_ net1015 VPWR _1584_ VGND net1228 net1005 sg13g2_o21ai_1
XFILLER_43_628 VPWR VGND sg13g2_decap_4
XFILLER_23_341 VPWR VGND sg13g2_decap_8
XFILLER_24_842 VPWR VGND sg13g2_fill_1
XFILLER_24_875 VPWR VGND sg13g2_decap_8
XFILLER_3_768 VPWR VGND sg13g2_decap_8
XFILLER_19_603 VPWR VGND sg13g2_decap_4
XFILLER_47_934 VPWR VGND sg13g2_decap_8
XFILLER_20_1018 VPWR VGND sg13g2_decap_8
XFILLER_33_138 VPWR VGND sg13g2_fill_2
XFILLER_15_875 VPWR VGND sg13g2_fill_1
XFILLER_30_801 VPWR VGND sg13g2_decap_8
X_3480_ _1901_ _1900_ net1267 _1886_ net1271 VPWR VGND sg13g2_a22oi_1
X_6173__99 VPWR VGND net99 sg13g2_tiehi
X_5150_ _0843_ net1127 _0842_ VPWR VGND sg13g2_nand2b_1
X_4101_ VPWR _2460_ net1181 VGND sg13g2_inv_1
X_5081_ VGND VPWR net1112 net471 _0781_ _0780_ sg13g2_a21oi_1
X_4032_ net1218 _2399_ _2400_ _2401_ VPWR VGND sg13g2_nor3_1
XFILLER_49_282 VPWR VGND sg13g2_fill_2
XFILLER_38_989 VPWR VGND sg13g2_decap_8
X_5983_ net32 VGND VPWR _0033_ s0.data_out\[19\]\[6\] clknet_leaf_36_clk sg13g2_dfrbpq_2
XFILLER_24_105 VPWR VGND sg13g2_decap_8
X_4934_ VGND VPWR _0643_ _0646_ _0649_ _0648_ sg13g2_a21oi_1
XFILLER_21_823 VPWR VGND sg13g2_fill_1
XFILLER_33_661 VPWR VGND sg13g2_decap_8
X_4865_ VPWR _0069_ net547 VGND sg13g2_inv_1
XFILLER_32_171 VPWR VGND sg13g2_decap_4
X_3816_ _2205_ net930 _2204_ VPWR VGND sg13g2_nand2_1
X_4796_ VGND VPWR _0522_ _0523_ _0059_ _0524_ sg13g2_a21oi_1
X_3747_ _2144_ _2143_ net1240 _2139_ net1233 VPWR VGND sg13g2_a22oi_1
X_3678_ _2080_ VPWR _2081_ VGND net1307 net420 sg13g2_o21ai_1
XFILLER_0_705 VPWR VGND sg13g2_decap_8
X_5417_ VGND VPWR net1105 _1085_ _1086_ _1056_ sg13g2_a21oi_1
X_5348_ VGND VPWR net1088 s0.data_out\[11\]\[2\] _1023_ _1022_ sg13g2_a21oi_1
X_5279_ _0959_ net1100 _0911_ _0960_ VPWR VGND sg13g2_a21o_1
XFILLER_29_923 VPWR VGND sg13g2_fill_2
X_6166__106 VPWR VGND net106 sg13g2_tiehi
XFILLER_44_948 VPWR VGND sg13g2_decap_8
XFILLER_28_477 VPWR VGND sg13g2_fill_2
XFILLER_8_816 VPWR VGND sg13g2_fill_1
XFILLER_23_193 VPWR VGND sg13g2_fill_2
XFILLER_7_29 VPWR VGND sg13g2_fill_1
XFILLER_7_359 VPWR VGND sg13g2_decap_4
XFILLER_2_0 VPWR VGND sg13g2_fill_1
Xfanout1322 net1323 net1322 VPWR VGND sg13g2_buf_8
Xfanout1300 net1350 net1300 VPWR VGND sg13g2_buf_8
Xfanout1311 net1312 net1311 VPWR VGND sg13g2_buf_8
Xfanout1333 net1339 net1333 VPWR VGND sg13g2_buf_8
Xfanout1344 net1347 net1344 VPWR VGND sg13g2_buf_8
XFILLER_47_731 VPWR VGND sg13g2_decap_8
XFILLER_4_1012 VPWR VGND sg13g2_decap_8
XFILLER_19_422 VPWR VGND sg13g2_decap_8
XFILLER_19_433 VPWR VGND sg13g2_fill_2
X_4650_ VGND VPWR _0391_ _0384_ net1233 sg13g2_or2_1
X_3601_ _2010_ net980 _2009_ VPWR VGND sg13g2_nand2b_1
X_4581_ net1156 s0.data_out\[17\]\[3\] _0327_ VPWR VGND sg13g2_and2_1
X_3532_ _1945_ _1948_ net1308 _1949_ VPWR VGND sg13g2_nand3_1
X_3463_ s0.data_out\[5\]\[2\] s0.data_out\[4\]\[2\] net987 _1884_ VPWR VGND sg13g2_mux2_1
X_6182_ net89 VGND VPWR _0232_ s0.data_out\[3\]\[6\] clknet_leaf_11_clk sg13g2_dfrbpq_2
X_5202_ net1100 net1075 _0891_ VPWR VGND sg13g2_nor2b_1
X_3394_ VGND VPWR _1819_ _1822_ _1825_ _1824_ sg13g2_a21oi_1
X_5133_ VPWR _0094_ net578 VGND sg13g2_inv_1
XFILLER_35_0 VPWR VGND sg13g2_decap_8
X_5064_ net1114 _0762_ _0767_ VPWR VGND sg13g2_nor2_1
X_4015_ _2388_ net1247 _2387_ VPWR VGND sg13g2_nand2_1
XFILLER_26_926 VPWR VGND sg13g2_decap_4
XFILLER_26_948 VPWR VGND sg13g2_fill_2
X_5966_ net50 VGND VPWR _0016_ s0.data_out\[20\]\[1\] clknet_leaf_37_clk sg13g2_dfrbpq_2
XFILLER_13_609 VPWR VGND sg13g2_fill_2
XFILLER_34_970 VPWR VGND sg13g2_decap_8
X_5897_ net1016 net1056 _1514_ VPWR VGND sg13g2_nor2b_1
X_4917_ _0621_ _0630_ _0632_ _0633_ _0634_ VPWR VGND sg13g2_nor4_1
X_4848_ _0568_ VPWR _0569_ VGND net1306 net416 sg13g2_o21ai_1
XFILLER_32_15 VPWR VGND sg13g2_decap_4
X_4779_ _0505_ _0506_ _0504_ _0508_ VPWR VGND sg13g2_nand3_1
XFILLER_10_1017 VPWR VGND sg13g2_decap_8
XFILLER_10_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_502 VPWR VGND sg13g2_decap_8
XFILLER_48_506 VPWR VGND sg13g2_decap_8
XFILLER_0_579 VPWR VGND sg13g2_decap_8
XFILLER_29_731 VPWR VGND sg13g2_fill_1
X_6033__250 VPWR VGND net250 sg13g2_tiehi
XFILLER_16_436 VPWR VGND sg13g2_fill_1
XFILLER_43_277 VPWR VGND sg13g2_decap_4
XFILLER_25_992 VPWR VGND sg13g2_decap_8
XFILLER_40_973 VPWR VGND sg13g2_decap_8
XFILLER_4_830 VPWR VGND sg13g2_decap_8
XFILLER_39_517 VPWR VGND sg13g2_fill_1
Xfanout1130 net1133 net1130 VPWR VGND sg13g2_buf_8
Xfanout1141 net1143 net1141 VPWR VGND sg13g2_buf_8
Xfanout1174 net1177 net1174 VPWR VGND sg13g2_buf_8
Xfanout1163 net1166 net1163 VPWR VGND sg13g2_buf_8
Xfanout1152 net1154 net1152 VPWR VGND sg13g2_buf_8
Xfanout1185 s0.shift_out\[19\][0] net1185 VPWR VGND sg13g2_buf_2
Xfanout1196 net333 net1196 VPWR VGND sg13g2_buf_8
XFILLER_19_230 VPWR VGND sg13g2_fill_2
XFILLER_19_285 VPWR VGND sg13g2_decap_8
XFILLER_23_907 VPWR VGND sg13g2_fill_2
X_5820_ net1243 _1443_ _1446_ VPWR VGND sg13g2_nor2_1
X_5751_ net1030 net1063 _1382_ VPWR VGND sg13g2_nor2b_1
XFILLER_34_277 VPWR VGND sg13g2_decap_8
XFILLER_34_299 VPWR VGND sg13g2_fill_1
X_4702_ net1145 net1065 _0437_ VPWR VGND sg13g2_nor2b_1
X_5682_ _1324_ _1326_ _1327_ VPWR VGND sg13g2_nor2_1
X_4633_ _0374_ net1164 s0.data_out\[17\]\[3\] VPWR VGND sg13g2_nand2_1
X_4564_ VGND VPWR _2808_ _0311_ _0312_ net1169 sg13g2_a21oi_1
X_3515_ net985 VPWR _1934_ VGND net1226 net974 sg13g2_o21ai_1
XFILLER_7_690 VPWR VGND sg13g2_fill_1
X_4495_ _2811_ net1181 _2810_ VPWR VGND sg13g2_nand2b_1
X_3446_ _1869_ net511 net998 VPWR VGND sg13g2_nand2b_1
X_3377_ _1798_ _1803_ _1809_ _1810_ VPWR VGND sg13g2_nor3_1
X_6165_ net107 VGND VPWR _0215_ s0.data_out\[4\]\[1\] clknet_leaf_5_clk sg13g2_dfrbpq_2
X_5116_ _0811_ VPWR _0812_ VGND _0807_ _0810_ sg13g2_o21ai_1
X_6017__267 VPWR VGND net267 sg13g2_tiehi
X_6096_ net182 VGND VPWR _0146_ s0.data_new_delayed\[2\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_5047_ net1264 _0726_ _0752_ VPWR VGND sg13g2_nor2_1
XFILLER_38_572 VPWR VGND sg13g2_fill_1
XFILLER_27_59 VPWR VGND sg13g2_fill_2
XFILLER_26_734 VPWR VGND sg13g2_fill_2
XFILLER_26_756 VPWR VGND sg13g2_fill_1
X_6163__109 VPWR VGND net109 sg13g2_tiehi
XFILLER_26_778 VPWR VGND sg13g2_decap_4
XFILLER_40_214 VPWR VGND sg13g2_decap_8
X_5949_ _1562_ _1560_ _1563_ VPWR VGND _1561_ sg13g2_nand3b_1
XFILLER_49_1024 VPWR VGND sg13g2_decap_4
XFILLER_4_126 VPWR VGND sg13g2_fill_2
XFILLER_4_159 VPWR VGND sg13g2_fill_1
XFILLER_1_844 VPWR VGND sg13g2_decap_8
XFILLER_0_343 VPWR VGND sg13g2_fill_2
XFILLER_29_561 VPWR VGND sg13g2_decap_4
XFILLER_1_1026 VPWR VGND sg13g2_fill_2
XFILLER_17_767 VPWR VGND sg13g2_decap_8
XFILLER_17_778 VPWR VGND sg13g2_fill_1
XFILLER_13_984 VPWR VGND sg13g2_decap_8
XFILLER_9_999 VPWR VGND sg13g2_decap_8
XFILLER_4_671 VPWR VGND sg13g2_fill_2
X_3300_ _1734_ _1737_ net1324 _1738_ VPWR VGND sg13g2_nand3_1
X_4280_ _2507_ _2617_ _2619_ _2620_ VPWR VGND sg13g2_nor3_1
X_3231_ VGND VPWR net1015 _1675_ _1676_ _1630_ sg13g2_a21oi_1
XFILLER_39_325 VPWR VGND sg13g2_decap_8
XFILLER_39_314 VPWR VGND sg13g2_fill_1
X_3162_ _1609_ _1612_ net1327 _1613_ VPWR VGND sg13g2_nand3_1
XFILLER_39_336 VPWR VGND sg13g2_fill_1
XFILLER_48_892 VPWR VGND sg13g2_decap_8
XFILLER_23_737 VPWR VGND sg13g2_fill_1
X_5803_ s0.data_out\[9\]\[3\] s0.data_out\[8\]\[3\] net1034 _1429_ VPWR VGND sg13g2_mux2_1
X_3995_ _2360_ _2366_ _2367_ _2368_ VPWR VGND sg13g2_or3_1
X_5734_ net1030 s0.data_out\[8\]\[1\] _1367_ VPWR VGND sg13g2_and2_1
X_5665_ _1310_ net1079 _1309_ VPWR VGND sg13g2_nand2b_1
XFILLER_31_792 VPWR VGND sg13g2_fill_1
X_4616_ VGND VPWR _0358_ net579 net1302 sg13g2_or2_1
X_5596_ net1036 s0.data_out\[9\]\[1\] _1248_ VPWR VGND sg13g2_and2_1
XFILLER_2_608 VPWR VGND sg13g2_decap_8
X_4547_ _0297_ VPWR _0298_ VGND net1171 _2740_ sg13g2_o21ai_1
X_4478_ _2795_ VPWR _2796_ VGND _2791_ _2794_ sg13g2_o21ai_1
X_6217_ net123 VGND VPWR _0267_ s0.data_out\[0\]\[5\] clknet_leaf_9_clk sg13g2_dfrbpq_2
Xfanout934 _2454_ net934 VPWR VGND sg13g2_buf_8
Xfanout912 net913 net912 VPWR VGND sg13g2_buf_8
Xfanout923 _2463_ net923 VPWR VGND sg13g2_buf_1
X_3429_ VPWR _0205_ _1854_ VGND sg13g2_inv_1
Xfanout945 net354 net945 VPWR VGND sg13g2_buf_8
Xfanout956 net958 net956 VPWR VGND sg13g2_buf_8
Xfanout967 net968 net967 VPWR VGND sg13g2_buf_1
X_6148_ net126 VGND VPWR _0198_ s0.shift_out\[6\][0] clknet_leaf_16_clk sg13g2_dfrbpq_1
Xfanout978 net979 net978 VPWR VGND sg13g2_buf_1
Xfanout989 s0.valid_out\[4\][0] net989 VPWR VGND sg13g2_buf_8
X_6079_ net200 VGND VPWR _0129_ s0.data_out\[11\]\[6\] clknet_leaf_20_clk sg13g2_dfrbpq_2
X_6030__253 VPWR VGND net253 sg13g2_tiehi
XFILLER_9_218 VPWR VGND sg13g2_decap_4
XFILLER_10_954 VPWR VGND sg13g2_decap_8
XFILLER_6_947 VPWR VGND sg13g2_decap_8
XFILLER_5_435 VPWR VGND sg13g2_fill_1
XFILLER_1_641 VPWR VGND sg13g2_decap_8
XFILLER_0_151 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_4
XFILLER_49_667 VPWR VGND sg13g2_decap_8
XFILLER_23_1027 VPWR VGND sg13g2_fill_2
XFILLER_36_317 VPWR VGND sg13g2_decap_4
XFILLER_17_520 VPWR VGND sg13g2_decap_8
XFILLER_28_91 VPWR VGND sg13g2_fill_2
XFILLER_45_851 VPWR VGND sg13g2_decap_8
X_3780_ net1299 VPWR _2175_ VGND net393 _2170_ sg13g2_o21ai_1
XFILLER_8_251 VPWR VGND sg13g2_fill_2
X_5450_ _1115_ _1116_ _1117_ VPWR VGND sg13g2_nor2_1
XFILLER_30_1009 VPWR VGND sg13g2_decap_8
X_4401_ VGND VPWR _2669_ _2727_ _2729_ net1246 sg13g2_a21oi_1
X_5381_ net1336 VPWR _1052_ VGND net938 _1051_ sg13g2_o21ai_1
XFILLER_5_73 VPWR VGND sg13g2_decap_8
X_4332_ net1182 net1057 _2664_ VPWR VGND sg13g2_nor2b_1
X_4263_ s0.data_out\[21\]\[4\] s0.data_out\[20\]\[4\] net1200 _2603_ VPWR VGND sg13g2_mux2_1
X_6002_ net283 VGND VPWR _0052_ s0.data_out\[17\]\[1\] clknet_leaf_35_clk sg13g2_dfrbpq_2
X_3214_ s0.data_out\[7\]\[0\] s0.data_out\[6\]\[0\] net1011 _1659_ VPWR VGND sg13g2_mux2_1
X_4194_ net1206 s0.data_out\[20\]\[3\] _2539_ VPWR VGND sg13g2_nor2_1
X_3145_ net1012 VPWR _1598_ VGND _1596_ _1597_ sg13g2_o21ai_1
XFILLER_23_501 VPWR VGND sg13g2_decap_8
XFILLER_10_206 VPWR VGND sg13g2_fill_1
XFILLER_23_567 VPWR VGND sg13g2_fill_1
X_3978_ s0.data_out\[1\]\[1\] s0.data_out\[0\]\[1\] net948 _2351_ VPWR VGND sg13g2_mux2_1
X_5717_ VGND VPWR _1353_ net1033 net398 sg13g2_or2_1
XFILLER_40_26 VPWR VGND sg13g2_decap_4
X_5648_ _1293_ VPWR _1294_ VGND _1289_ _1292_ sg13g2_o21ai_1
X_5579_ VGND VPWR _1234_ net1043 s0.was_valid_out\[9\][0] sg13g2_or2_1
XFILLER_2_438 VPWR VGND sg13g2_decap_8
Xhold262 s0.data_out\[18\]\[6\] VPWR VGND net558 sg13g2_dlygate4sd3_1
Xhold251 _0583_ VPWR VGND net547 sg13g2_dlygate4sd3_1
Xhold240 s0.data_out\[11\]\[1\] VPWR VGND net536 sg13g2_dlygate4sd3_1
XFILLER_49_35 VPWR VGND sg13g2_decap_8
Xhold273 s0.data_out\[5\]\[7\] VPWR VGND net569 sg13g2_dlygate4sd3_1
XFILLER_46_1027 VPWR VGND sg13g2_fill_2
Xhold284 _0359_ VPWR VGND net580 sg13g2_dlygate4sd3_1
Xhold295 s0.data_out\[16\]\[7\] VPWR VGND net591 sg13g2_dlygate4sd3_1
XFILLER_18_317 VPWR VGND sg13g2_fill_1
XFILLER_46_648 VPWR VGND sg13g2_decap_4
XFILLER_27_851 VPWR VGND sg13g2_decap_8
XFILLER_14_501 VPWR VGND sg13g2_decap_8
XFILLER_26_394 VPWR VGND sg13g2_fill_2
XFILLER_42_887 VPWR VGND sg13g2_decap_8
XFILLER_6_711 VPWR VGND sg13g2_decap_8
X_6185__86 VPWR VGND net86 sg13g2_tiehi
XFILLER_5_221 VPWR VGND sg13g2_fill_1
XFILLER_5_232 VPWR VGND sg13g2_decap_8
XFILLER_2_994 VPWR VGND sg13g2_decap_8
XFILLER_49_464 VPWR VGND sg13g2_decap_8
XFILLER_36_158 VPWR VGND sg13g2_fill_2
X_4950_ net1138 VPWR _0662_ VGND _0660_ _0661_ sg13g2_o21ai_1
X_3901_ VGND VPWR net1222 net947 _2284_ _2283_ sg13g2_a21oi_1
X_4881_ VGND VPWR _0543_ _0596_ _0598_ net1277 sg13g2_a21oi_1
X_3832_ VGND VPWR _2140_ _2218_ _2219_ net964 sg13g2_a21oi_1
X_5502_ net1080 net1055 _1162_ VPWR VGND sg13g2_nor2b_1
X_3763_ _2158_ VPWR _2160_ VGND _2130_ _2135_ sg13g2_o21ai_1
X_3694_ _2094_ VPWR _2095_ VGND net1307 net441 sg13g2_o21ai_1
X_5433_ _1101_ net1091 _1043_ _1102_ VPWR VGND sg13g2_a21o_1
X_5364_ VGND VPWR net1092 net330 _1037_ _1036_ sg13g2_a21oi_1
X_4315_ net1178 net1065 _2649_ VPWR VGND sg13g2_nor2b_1
X_5295_ VGND VPWR _0976_ _0968_ net1236 sg13g2_or2_1
X_4246_ _2585_ net1191 _2536_ _2586_ VPWR VGND sg13g2_a21o_1
X_4177_ VGND VPWR net1206 _2481_ _2524_ net1202 sg13g2_a21oi_1
XFILLER_28_604 VPWR VGND sg13g2_fill_2
X_3128_ net1326 net313 _0175_ VPWR VGND sg13g2_and2_1
XFILLER_24_821 VPWR VGND sg13g2_fill_1
XFILLER_24_887 VPWR VGND sg13g2_decap_4
XFILLER_13_1026 VPWR VGND sg13g2_fill_2
X_6182__89 VPWR VGND net89 sg13g2_tiehi
XFILLER_4_4 VPWR VGND sg13g2_decap_4
XFILLER_3_747 VPWR VGND sg13g2_decap_8
XFILLER_47_913 VPWR VGND sg13g2_decap_8
XFILLER_46_412 VPWR VGND sg13g2_fill_2
XFILLER_18_114 VPWR VGND sg13g2_fill_1
XFILLER_27_670 VPWR VGND sg13g2_fill_1
XFILLER_14_364 VPWR VGND sg13g2_decap_8
XFILLER_41_91 VPWR VGND sg13g2_fill_1
XFILLER_10_592 VPWR VGND sg13g2_fill_2
XFILLER_6_585 VPWR VGND sg13g2_fill_2
X_4100_ VPWR _2459_ net952 VGND sg13g2_inv_1
X_5080_ net1112 net1070 _0780_ VPWR VGND sg13g2_nor2b_1
XFILLER_2_791 VPWR VGND sg13g2_decap_8
X_4031_ net1073 net940 _2400_ VPWR VGND sg13g2_nor2b_1
XFILLER_38_968 VPWR VGND sg13g2_decap_8
X_5982_ net33 VGND VPWR _0032_ s0.data_out\[19\]\[5\] clknet_leaf_3_clk sg13g2_dfrbpq_2
X_4933_ _0647_ VPWR _0648_ VGND net1125 _0641_ sg13g2_o21ai_1
XFILLER_36_1015 VPWR VGND sg13g2_decap_8
X_4864_ _0582_ VPWR _0583_ VGND _0578_ _0581_ sg13g2_o21ai_1
X_3815_ s0.data_out\[1\]\[4\] s0.data_out\[2\]\[4\] net966 _2204_ VPWR VGND sg13g2_mux2_1
X_4795_ VGND VPWR _0524_ net1208 net308 sg13g2_or2_1
XFILLER_20_345 VPWR VGND sg13g2_fill_1
X_3746_ VGND VPWR net973 _2142_ _2143_ _2104_ sg13g2_a21oi_1
X_6159__114 VPWR VGND net114 sg13g2_tiehi
X_5416_ _1084_ net1091 _1057_ _1085_ VPWR VGND sg13g2_a21o_1
X_3677_ _2076_ _2079_ net1307 _2080_ VPWR VGND sg13g2_nand3_1
X_5347_ net1089 net1066 _1022_ VPWR VGND sg13g2_nor2b_1
X_5278_ s0.data_out\[13\]\[3\] s0.data_out\[12\]\[3\] net1108 _0959_ VPWR VGND sg13g2_mux2_1
X_4229_ _0010_ _2565_ _2569_ _2472_ net1216 VPWR VGND sg13g2_a22oi_1
XFILLER_29_957 VPWR VGND sg13g2_fill_1
XFILLER_44_927 VPWR VGND sg13g2_decap_8
XFILLER_43_459 VPWR VGND sg13g2_fill_1
XFILLER_43_448 VPWR VGND sg13g2_decap_8
XFILLER_11_356 VPWR VGND sg13g2_decap_8
XFILLER_7_327 VPWR VGND sg13g2_decap_4
XFILLER_11_50 VPWR VGND sg13g2_decap_8
Xfanout1301 net1302 net1301 VPWR VGND sg13g2_buf_8
Xfanout1323 net1349 net1323 VPWR VGND sg13g2_buf_8
Xfanout1312 net1315 net1312 VPWR VGND sg13g2_buf_8
Xfanout1334 net1335 net1334 VPWR VGND sg13g2_buf_8
Xfanout1345 net1347 net1345 VPWR VGND sg13g2_buf_1
XFILLER_47_710 VPWR VGND sg13g2_decap_8
XFILLER_47_787 VPWR VGND sg13g2_decap_8
XFILLER_43_982 VPWR VGND sg13g2_decap_8
XFILLER_42_481 VPWR VGND sg13g2_fill_2
XFILLER_14_183 VPWR VGND sg13g2_fill_2
X_4580_ _0326_ net925 _0325_ VPWR VGND sg13g2_nand2_1
X_3600_ VGND VPWR net969 _2008_ _2009_ _1947_ sg13g2_a21oi_1
X_3531_ net980 VPWR _1948_ VGND _1946_ _1947_ sg13g2_o21ai_1
X_3462_ _1883_ net987 net533 VPWR VGND sg13g2_nand2_1
X_6181_ net90 VGND VPWR _0231_ s0.data_out\[3\]\[5\] clknet_leaf_11_clk sg13g2_dfrbpq_2
X_3393_ _1823_ VPWR _1824_ VGND net985 _1817_ sg13g2_o21ai_1
X_5201_ net1100 s0.data_out\[12\]\[0\] _0890_ VPWR VGND sg13g2_and2_1
X_5132_ _0825_ VPWR _0826_ VGND _0821_ _0824_ sg13g2_o21ai_1
X_5063_ _0763_ VPWR _0766_ VGND net346 net1119 sg13g2_o21ai_1
X_4014_ _2327_ _2386_ _2387_ VPWR VGND sg13g2_and2_1
XFILLER_37_242 VPWR VGND sg13g2_fill_2
XFILLER_38_787 VPWR VGND sg13g2_decap_8
XFILLER_16_17 VPWR VGND sg13g2_fill_2
XFILLER_25_448 VPWR VGND sg13g2_fill_1
XFILLER_41_919 VPWR VGND sg13g2_decap_8
X_5965_ net51 VGND VPWR _0015_ s0.data_out\[20\]\[0\] clknet_leaf_37_clk sg13g2_dfrbpq_2
X_5896_ VGND VPWR _1450_ _1512_ _1513_ net1025 sg13g2_a21oi_1
X_4916_ _0633_ _0631_ _0625_ VPWR VGND sg13g2_nand2b_1
XFILLER_21_621 VPWR VGND sg13g2_decap_4
X_4847_ _0564_ _0567_ net1319 _0568_ VPWR VGND sg13g2_nand3_1
XFILLER_20_131 VPWR VGND sg13g2_decap_8
XFILLER_20_175 VPWR VGND sg13g2_decap_8
X_4778_ _0507_ _0504_ _0505_ _0506_ VPWR VGND sg13g2_and3_1
X_3729_ VGND VPWR net959 _2125_ _2126_ _2064_ sg13g2_a21oi_1
X_6172__100 VPWR VGND net100 sg13g2_tiehi
XFILLER_0_558 VPWR VGND sg13g2_decap_8
XFILLER_44_724 VPWR VGND sg13g2_fill_1
XFILLER_17_927 VPWR VGND sg13g2_decap_8
XFILLER_29_776 VPWR VGND sg13g2_fill_2
XFILLER_43_223 VPWR VGND sg13g2_fill_2
XFILLER_43_267 VPWR VGND sg13g2_fill_2
XFILLER_40_952 VPWR VGND sg13g2_decap_8
XFILLER_12_676 VPWR VGND sg13g2_fill_2
XFILLER_4_886 VPWR VGND sg13g2_decap_8
Xfanout1131 net1133 net1131 VPWR VGND sg13g2_buf_8
Xfanout1120 s0.valid_out\[13\][0] net1120 VPWR VGND sg13g2_buf_8
Xfanout1164 net1166 net1164 VPWR VGND sg13g2_buf_8
Xfanout1142 net1143 net1142 VPWR VGND sg13g2_buf_8
Xfanout1153 net1154 net1153 VPWR VGND sg13g2_buf_2
Xfanout1186 net1189 net1186 VPWR VGND sg13g2_buf_8
Xfanout1175 net1177 net1175 VPWR VGND sg13g2_buf_1
Xfanout1197 net333 net1197 VPWR VGND sg13g2_buf_1
XFILLER_47_595 VPWR VGND sg13g2_decap_8
XFILLER_19_297 VPWR VGND sg13g2_decap_4
XFILLER_34_256 VPWR VGND sg13g2_decap_8
XFILLER_16_993 VPWR VGND sg13g2_decap_8
XFILLER_22_418 VPWR VGND sg13g2_decap_4
XFILLER_22_429 VPWR VGND sg13g2_fill_1
X_5750_ net1030 s0.data_out\[8\]\[3\] _1381_ VPWR VGND sg13g2_and2_1
X_4701_ VGND VPWR _0360_ _0435_ _0436_ net1161 sg13g2_a21oi_1
X_5681_ _1326_ _1322_ _1325_ VPWR VGND sg13g2_nand2_1
X_4632_ VPWR VGND _0305_ net1281 _0371_ net1275 _0373_ _0368_ sg13g2_a221oi_1
XFILLER_30_473 VPWR VGND sg13g2_fill_2
XFILLER_31_985 VPWR VGND sg13g2_decap_8
XFILLER_33_1018 VPWR VGND sg13g2_decap_8
XFILLER_8_84 VPWR VGND sg13g2_decap_8
X_4563_ _0311_ s0.data_out\[17\]\[1\] net1175 VPWR VGND sg13g2_nand2b_1
X_3514_ net1310 net317 _0211_ VPWR VGND sg13g2_and2_1
X_4494_ VGND VPWR net1168 _2809_ _2810_ _2758_ sg13g2_a21oi_1
X_6156__117 VPWR VGND net117 sg13g2_tiehi
X_3445_ VPWR _0207_ _1868_ VGND sg13g2_inv_1
X_6164_ net108 VGND VPWR _0214_ s0.data_out\[4\]\[0\] clknet_leaf_4_clk sg13g2_dfrbpq_2
X_3376_ net1250 _1801_ _1809_ VPWR VGND sg13g2_nor2_1
X_5115_ VGND VPWR _0811_ net548 net1322 sg13g2_or2_1
X_6095_ net183 VGND VPWR _0145_ s0.data_new_delayed\[1\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_5046_ _0687_ _0750_ net1250 _0751_ VPWR VGND sg13g2_nand3_1
XFILLER_26_713 VPWR VGND sg13g2_decap_4
XFILLER_14_908 VPWR VGND sg13g2_decap_4
XFILLER_25_234 VPWR VGND sg13g2_fill_2
XFILLER_25_245 VPWR VGND sg13g2_decap_8
X_5948_ VGND VPWR _1562_ _1555_ net1237 sg13g2_or2_1
XFILLER_43_59 VPWR VGND sg13g2_fill_2
XFILLER_21_451 VPWR VGND sg13g2_decap_8
XFILLER_21_462 VPWR VGND sg13g2_fill_2
XFILLER_22_985 VPWR VGND sg13g2_decap_8
X_5879_ s0.data_out\[7\]\[3\] s0.data_out\[8\]\[3\] net1031 _1498_ VPWR VGND sg13g2_mux2_1
XFILLER_5_606 VPWR VGND sg13g2_decap_4
XFILLER_49_1003 VPWR VGND sg13g2_decap_8
XFILLER_4_116 VPWR VGND sg13g2_fill_2
XFILLER_1_823 VPWR VGND sg13g2_decap_8
XFILLER_0_322 VPWR VGND sg13g2_decap_8
XFILLER_49_849 VPWR VGND sg13g2_decap_8
XFILLER_29_540 VPWR VGND sg13g2_fill_1
XFILLER_1_1005 VPWR VGND sg13g2_decap_8
XFILLER_29_584 VPWR VGND sg13g2_decap_8
XFILLER_17_82 VPWR VGND sg13g2_decap_8
XFILLER_44_587 VPWR VGND sg13g2_fill_2
XFILLER_16_289 VPWR VGND sg13g2_decap_4
XFILLER_13_963 VPWR VGND sg13g2_decap_8
XFILLER_9_978 VPWR VGND sg13g2_decap_8
X_3230_ _1674_ net1005 _1631_ _1675_ VPWR VGND sg13g2_a21o_1
X_3161_ net1012 VPWR _1612_ VGND _1610_ _1611_ sg13g2_o21ai_1
XFILLER_48_871 VPWR VGND sg13g2_decap_8
X_5802_ VPWR VGND _1426_ _1427_ _1422_ net1213 _1428_ _1417_ sg13g2_a221oi_1
X_3994_ net1211 _2350_ _2367_ VPWR VGND sg13g2_nor2_1
XFILLER_13_29 VPWR VGND sg13g2_fill_1
X_5733_ _1366_ net919 _1365_ VPWR VGND sg13g2_nand2_1
X_5664_ VGND VPWR net1036 _1308_ _1309_ _1263_ sg13g2_a21oi_1
X_4615_ net1301 VPWR _0357_ VGND net925 _0356_ sg13g2_o21ai_1
X_6023__261 VPWR VGND net261 sg13g2_tiehi
X_5595_ _1247_ net934 _1246_ VPWR VGND sg13g2_nand2_1
X_4546_ VPWR _0297_ _0296_ VGND sg13g2_inv_1
X_4477_ VGND VPWR _2795_ net551 net1288 sg13g2_or2_1
Xfanout924 _2462_ net924 VPWR VGND sg13g2_buf_8
Xfanout913 _2494_ net913 VPWR VGND sg13g2_buf_8
X_3428_ _1853_ VPWR _1854_ VGND net1311 net415 sg13g2_o21ai_1
X_6216_ net136 VGND VPWR _0266_ s0.data_out\[0\]\[4\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_6147_ net127 VGND VPWR _0197_ s0.data_out\[6\]\[7\] clknet_leaf_17_clk sg13g2_dfrbpq_2
Xfanout957 net958 net957 VPWR VGND sg13g2_buf_2
X_3359_ s0.data_out\[6\]\[6\] s0.data_out\[5\]\[6\] net999 _1792_ VPWR VGND sg13g2_mux2_1
Xfanout968 s0.valid_out\[2\][0] net968 VPWR VGND sg13g2_buf_8
Xfanout935 _2453_ net935 VPWR VGND sg13g2_buf_8
Xfanout946 net948 net946 VPWR VGND sg13g2_buf_8
Xfanout979 s0.valid_out\[3\][0] net979 VPWR VGND sg13g2_buf_8
X_6078_ net201 VGND VPWR _0128_ s0.data_out\[11\]\[5\] clknet_leaf_26_clk sg13g2_dfrbpq_2
XFILLER_39_882 VPWR VGND sg13g2_fill_2
X_5029_ s0.data_out\[15\]\[6\] s0.data_out\[14\]\[6\] net1130 _0734_ VPWR VGND sg13g2_mux2_1
XFILLER_14_727 VPWR VGND sg13g2_fill_2
XFILLER_10_933 VPWR VGND sg13g2_decap_8
X_6197__73 VPWR VGND net73 sg13g2_tiehi
XFILLER_22_782 VPWR VGND sg13g2_fill_2
XFILLER_6_926 VPWR VGND sg13g2_decap_8
XFILLER_1_620 VPWR VGND sg13g2_decap_8
XFILLER_49_646 VPWR VGND sg13g2_decap_8
XFILLER_37_808 VPWR VGND sg13g2_fill_2
XFILLER_0_185 VPWR VGND sg13g2_decap_8
XFILLER_1_697 VPWR VGND sg13g2_decap_8
XFILLER_23_1006 VPWR VGND sg13g2_decap_8
XFILLER_45_830 VPWR VGND sg13g2_decap_8
XFILLER_29_381 VPWR VGND sg13g2_decap_8
XFILLER_17_554 VPWR VGND sg13g2_decap_8
XFILLER_8_230 VPWR VGND sg13g2_fill_2
X_6007__278 VPWR VGND net278 sg13g2_tiehi
X_4400_ _2669_ _2727_ net1246 _2728_ VPWR VGND sg13g2_nand3_1
X_5380_ VGND VPWR net1091 net527 _1051_ _1050_ sg13g2_a21oi_1
X_4331_ net1182 s0.data_out\[19\]\[4\] _2663_ VPWR VGND sg13g2_and2_1
X_4262_ _2601_ _2599_ _2602_ VPWR VGND _2600_ sg13g2_nand3b_1
X_6001_ net284 VGND VPWR _0051_ s0.data_out\[17\]\[0\] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_3213_ _1602_ _1657_ net1278 _1658_ VPWR VGND sg13g2_nand3_1
X_4193_ net366 net1206 _2538_ VPWR VGND sg13g2_nor2b_1
X_3144_ net1001 net1074 _1597_ VPWR VGND sg13g2_nor2b_1
XFILLER_24_17 VPWR VGND sg13g2_decap_4
XFILLER_11_719 VPWR VGND sg13g2_decap_8
X_3977_ _2306_ VPWR _2350_ VGND net928 _2349_ sg13g2_o21ai_1
X_5716_ _1351_ VPWR _1352_ VGND net1038 _1230_ sg13g2_o21ai_1
X_6194__76 VPWR VGND net76 sg13g2_tiehi
XFILLER_40_49 VPWR VGND sg13g2_decap_8
X_5647_ VGND VPWR _1293_ net531 net1346 sg13g2_or2_1
XFILLER_3_929 VPWR VGND sg13g2_decap_8
X_5578_ _1232_ VPWR _1233_ VGND net1082 _1116_ sg13g2_o21ai_1
XFILLER_46_1006 VPWR VGND sg13g2_decap_8
X_4529_ _2777_ _0281_ net1254 _0282_ VPWR VGND sg13g2_nand3_1
Xhold252 s0.data_out\[14\]\[5\] VPWR VGND net548 sg13g2_dlygate4sd3_1
X_6097__181 VPWR VGND net181 sg13g2_tiehi
Xhold241 s0.data_out\[6\]\[1\] VPWR VGND net537 sg13g2_dlygate4sd3_1
Xhold230 s0.data_out\[8\]\[1\] VPWR VGND net526 sg13g2_dlygate4sd3_1
XFILLER_49_14 VPWR VGND sg13g2_decap_8
Xhold263 _0352_ VPWR VGND net559 sg13g2_dlygate4sd3_1
Xhold296 s0.data_out\[20\]\[6\] VPWR VGND net592 sg13g2_dlygate4sd3_1
Xhold274 s0.data_out\[18\]\[5\] VPWR VGND net570 sg13g2_dlygate4sd3_1
Xhold285 s0.data_out\[5\]\[2\] VPWR VGND net581 sg13g2_dlygate4sd3_1
XFILLER_18_307 VPWR VGND sg13g2_decap_4
XFILLER_27_885 VPWR VGND sg13g2_decap_8
XFILLER_42_866 VPWR VGND sg13g2_decap_8
XFILLER_14_524 VPWR VGND sg13g2_fill_1
XFILLER_14_579 VPWR VGND sg13g2_decap_8
XFILLER_14_61 VPWR VGND sg13g2_decap_8
XFILLER_10_774 VPWR VGND sg13g2_decap_4
XFILLER_5_255 VPWR VGND sg13g2_decap_8
XFILLER_5_288 VPWR VGND sg13g2_decap_8
XFILLER_30_93 VPWR VGND sg13g2_decap_8
XFILLER_2_973 VPWR VGND sg13g2_decap_8
XFILLER_1_483 VPWR VGND sg13g2_decap_8
XFILLER_49_443 VPWR VGND sg13g2_decap_8
XFILLER_39_80 VPWR VGND sg13g2_decap_8
XFILLER_36_104 VPWR VGND sg13g2_fill_2
XFILLER_36_137 VPWR VGND sg13g2_fill_1
X_6013__271 VPWR VGND net271 sg13g2_tiehi
XFILLER_45_682 VPWR VGND sg13g2_decap_4
XFILLER_17_373 VPWR VGND sg13g2_decap_4
XFILLER_18_874 VPWR VGND sg13g2_decap_8
X_3900_ net952 VPWR _2283_ VGND net1225 net943 sg13g2_o21ai_1
X_4880_ _0543_ _0596_ net1277 _0597_ VPWR VGND sg13g2_nand3_1
XFILLER_33_833 VPWR VGND sg13g2_decap_8
X_3831_ _2218_ s0.data_out\[1\]\[6\] net966 VPWR VGND sg13g2_nand2b_1
X_3762_ _2155_ VPWR _2159_ VGND net1255 _2151_ sg13g2_o21ai_1
XFILLER_20_527 VPWR VGND sg13g2_fill_2
XFILLER_32_376 VPWR VGND sg13g2_decap_8
X_5501_ VGND VPWR _1100_ _1160_ _1161_ net1093 sg13g2_a21oi_1
X_3693_ _2090_ _2093_ net1307 _2094_ VPWR VGND sg13g2_nand3_1
X_5432_ s0.data_out\[12\]\[5\] s0.data_out\[11\]\[5\] net1098 _1101_ VPWR VGND sg13g2_mux2_1
X_6020__264 VPWR VGND net264 sg13g2_tiehi
X_5363_ net1092 net1059 _1036_ VPWR VGND sg13g2_nor2b_1
X_6191__79 VPWR VGND net79 sg13g2_tiehi
X_4314_ VGND VPWR _2570_ _2647_ _2648_ net1193 sg13g2_a21oi_1
X_5294_ net1236 _0968_ _0975_ VPWR VGND sg13g2_nor2_1
X_4245_ s0.data_out\[21\]\[3\] s0.data_out\[20\]\[3\] net1198 _2585_ VPWR VGND sg13g2_mux2_1
X_4176_ net1202 VPWR _2523_ VGND _2521_ _2522_ sg13g2_o21ai_1
X_3127_ VGND VPWR _1578_ _1582_ _0174_ _1583_ sg13g2_a21oi_1
XFILLER_28_638 VPWR VGND sg13g2_decap_8
XFILLER_23_365 VPWR VGND sg13g2_decap_8
XFILLER_11_516 VPWR VGND sg13g2_decap_4
XFILLER_13_1005 VPWR VGND sg13g2_decap_8
XFILLER_3_726 VPWR VGND sg13g2_decap_8
XFILLER_47_969 VPWR VGND sg13g2_decap_8
XFILLER_46_457 VPWR VGND sg13g2_decap_4
XFILLER_15_811 VPWR VGND sg13g2_decap_8
XFILLER_15_822 VPWR VGND sg13g2_fill_1
XFILLER_34_619 VPWR VGND sg13g2_fill_1
XFILLER_29_1023 VPWR VGND sg13g2_decap_4
X_6181__90 VPWR VGND net90 sg13g2_tiehi
XFILLER_2_770 VPWR VGND sg13g2_decap_8
XFILLER_38_914 VPWR VGND sg13g2_fill_1
X_4030_ VGND VPWR net946 net377 _2399_ net940 sg13g2_a21oi_1
XFILLER_38_947 VPWR VGND sg13g2_decap_8
XFILLER_37_446 VPWR VGND sg13g2_fill_1
XFILLER_2_97 VPWR VGND sg13g2_fill_2
X_5981_ net34 VGND VPWR _0031_ s0.data_out\[19\]\[4\] clknet_leaf_3_clk sg13g2_dfrbpq_2
X_4932_ net921 VPWR _0647_ VGND net378 net1143 sg13g2_o21ai_1
XFILLER_33_630 VPWR VGND sg13g2_fill_2
X_6087__191 VPWR VGND net191 sg13g2_tiehi
X_4863_ VGND VPWR _0582_ net546 net1318 sg13g2_or2_1
X_4794_ VPWR VGND _0507_ _0419_ _0521_ _0495_ _0523_ _0519_ sg13g2_a221oi_1
X_3814_ VPWR _0241_ net447 VGND sg13g2_inv_1
X_3745_ _2141_ net964 _2105_ _2142_ VPWR VGND sg13g2_a21o_1
X_5415_ s0.data_out\[12\]\[7\] s0.data_out\[11\]\[7\] net1098 _1084_ VPWR VGND sg13g2_mux2_1
X_3676_ net971 VPWR _2079_ VGND _2077_ _2078_ sg13g2_o21ai_1
X_5346_ VGND VPWR _0944_ _1020_ _1021_ net1102 sg13g2_a21oi_1
X_5277_ VPWR VGND _0956_ _0957_ _0952_ net1212 _0958_ _0947_ sg13g2_a221oi_1
X_6094__184 VPWR VGND net184 sg13g2_tiehi
X_4228_ net1216 _2568_ _2569_ VPWR VGND sg13g2_nor2_1
XFILLER_29_903 VPWR VGND sg13g2_fill_2
XFILLER_29_936 VPWR VGND sg13g2_fill_2
XFILLER_44_906 VPWR VGND sg13g2_decap_8
X_4159_ _2505_ _2508_ _2509_ VPWR VGND sg13g2_nor2_1
XFILLER_28_446 VPWR VGND sg13g2_decap_8
XFILLER_28_479 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_35_clk clknet_3_1__leaf_clk clknet_leaf_35_clk VPWR VGND sg13g2_buf_8
XFILLER_12_803 VPWR VGND sg13g2_decap_4
XFILLER_11_302 VPWR VGND sg13g2_fill_2
XFILLER_23_195 VPWR VGND sg13g2_fill_1
Xfanout1313 net1315 net1313 VPWR VGND sg13g2_buf_8
Xfanout1302 net1303 net1302 VPWR VGND sg13g2_buf_2
Xfanout1335 net1339 net1335 VPWR VGND sg13g2_buf_8
Xfanout1324 net1326 net1324 VPWR VGND sg13g2_buf_8
Xfanout1346 net1347 net1346 VPWR VGND sg13g2_buf_8
XFILLER_19_402 VPWR VGND sg13g2_decap_8
XFILLER_19_413 VPWR VGND sg13g2_fill_1
XFILLER_47_766 VPWR VGND sg13g2_decap_8
XFILLER_43_961 VPWR VGND sg13g2_decap_8
XFILLER_15_641 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_26_clk clknet_3_5__leaf_clk clknet_leaf_26_clk VPWR VGND sg13g2_buf_8
XFILLER_15_685 VPWR VGND sg13g2_decap_4
XFILLER_15_696 VPWR VGND sg13g2_decap_4
X_3530_ net969 net1076 _1947_ VPWR VGND sg13g2_nor2b_1
X_3461_ VPWR _0209_ _1882_ VGND sg13g2_inv_1
XFILLER_6_383 VPWR VGND sg13g2_fill_2
X_3392_ net915 VPWR _1823_ VGND net353 net998 sg13g2_o21ai_1
X_6180_ net91 VGND VPWR _0230_ s0.data_out\[3\]\[4\] clknet_leaf_14_clk sg13g2_dfrbpq_2
X_5200_ _0889_ net935 _0888_ VPWR VGND sg13g2_nand2_1
X_5131_ VGND VPWR _0825_ net577 net1333 sg13g2_or2_1
X_5062_ _0764_ VPWR _0765_ VGND net1126 _0642_ sg13g2_o21ai_1
XFILLER_42_1020 VPWR VGND sg13g2_decap_8
X_4013_ _2386_ net952 _2385_ VPWR VGND sg13g2_nand2b_1
XFILLER_37_221 VPWR VGND sg13g2_decap_8
XFILLER_19_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_17_clk clknet_3_6__leaf_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
X_5964_ net52 VGND VPWR _0014_ s0.valid_out\[20\][0] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_5895_ _1512_ s0.data_out\[7\]\[5\] net1032 VPWR VGND sg13g2_nand2b_1
X_4915_ _0626_ VPWR _0632_ VGND net1264 _0607_ sg13g2_o21ai_1
X_4846_ net1150 VPWR _0567_ VGND _0565_ _0566_ sg13g2_o21ai_1
XFILLER_21_633 VPWR VGND sg13g2_decap_8
XFILLER_20_165 VPWR VGND sg13g2_fill_1
X_4777_ VGND VPWR _0506_ _0499_ net1240 sg13g2_or2_1
X_3728_ s0.data_out\[3\]\[0\] s0.data_out\[2\]\[0\] net965 _2125_ VPWR VGND sg13g2_mux2_1
X_3659_ net959 net1076 _2064_ VPWR VGND sg13g2_nor2b_1
XFILLER_0_537 VPWR VGND sg13g2_decap_8
X_5329_ s0.data_out\[11\]\[0\] s0.data_out\[12\]\[0\] net1108 _1006_ VPWR VGND sg13g2_mux2_1
X_6213__175 VPWR VGND net175 sg13g2_tiehi
XFILLER_28_265 VPWR VGND sg13g2_decap_8
XFILLER_16_427 VPWR VGND sg13g2_decap_8
XFILLER_44_769 VPWR VGND sg13g2_decap_4
XFILLER_40_931 VPWR VGND sg13g2_decap_8
XFILLER_40_920 VPWR VGND sg13g2_fill_2
XFILLER_12_622 VPWR VGND sg13g2_fill_2
XFILLER_19_1022 VPWR VGND sg13g2_decap_8
XFILLER_8_626 VPWR VGND sg13g2_decap_4
XFILLER_7_114 VPWR VGND sg13g2_fill_2
XFILLER_11_143 VPWR VGND sg13g2_decap_4
XFILLER_4_865 VPWR VGND sg13g2_decap_8
XFILLER_3_342 VPWR VGND sg13g2_decap_8
Xfanout1121 s0.valid_out\[13\][0] net1121 VPWR VGND sg13g2_buf_8
Xfanout1110 net1111 net1110 VPWR VGND sg13g2_buf_8
Xfanout1132 net1133 net1132 VPWR VGND sg13g2_buf_2
XFILLER_26_1015 VPWR VGND sg13g2_decap_8
Xfanout1165 net1166 net1165 VPWR VGND sg13g2_buf_2
Xfanout1154 s0.valid_out\[16\][0] net1154 VPWR VGND sg13g2_buf_8
Xfanout1143 net601 net1143 VPWR VGND sg13g2_buf_8
Xfanout1198 net1201 net1198 VPWR VGND sg13g2_buf_8
Xfanout1187 net1189 net1187 VPWR VGND sg13g2_buf_1
Xfanout1176 net1177 net1176 VPWR VGND sg13g2_buf_8
XFILLER_19_232 VPWR VGND sg13g2_fill_1
XFILLER_47_585 VPWR VGND sg13g2_decap_4
X_6149__125 VPWR VGND net125 sg13g2_tiehi
XFILLER_16_961 VPWR VGND sg13g2_decap_8
XFILLER_23_909 VPWR VGND sg13g2_fill_1
X_4700_ _0435_ net422 net1164 VPWR VGND sg13g2_nand2b_1
XFILLER_31_942 VPWR VGND sg13g2_decap_4
XFILLER_31_964 VPWR VGND sg13g2_decap_8
X_6084__194 VPWR VGND net194 sg13g2_tiehi
X_5680_ VGND VPWR _1325_ _1317_ net1237 sg13g2_or2_1
X_4631_ _0364_ VPWR _0372_ VGND net1275 _0368_ sg13g2_o21ai_1
X_4562_ VPWR _0039_ _0310_ VGND sg13g2_inv_1
X_3513_ VGND VPWR _1928_ _1932_ _0210_ _1933_ sg13g2_a21oi_1
X_4493_ s0.data_out\[19\]\[1\] s0.data_out\[18\]\[1\] net1174 _2809_ VPWR VGND sg13g2_mux2_1
X_3444_ _1867_ VPWR _1868_ VGND net1314 net352 sg13g2_o21ai_1
Xclkbuf_leaf_6_clk clknet_3_2__leaf_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
XFILLER_40_0 VPWR VGND sg13g2_decap_8
X_6163_ net109 VGND VPWR _0213_ s0.valid_out\[4\][0] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_3375_ _1741_ _1806_ net1258 _1808_ VPWR VGND sg13g2_nand3_1
X_6091__187 VPWR VGND net187 sg13g2_tiehi
X_5114_ net1322 VPWR _0810_ VGND net937 _0809_ sg13g2_o21ai_1
X_6094_ net184 VGND VPWR _0144_ s0.data_new_delayed\[0\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_5045_ _0750_ net1139 _0749_ VPWR VGND sg13g2_nand2b_1
XFILLER_25_213 VPWR VGND sg13g2_decap_8
X_5947_ net1242 _1559_ _1561_ VPWR VGND sg13g2_nor2_1
XFILLER_22_920 VPWR VGND sg13g2_fill_2
XFILLER_40_227 VPWR VGND sg13g2_fill_1
XFILLER_22_942 VPWR VGND sg13g2_fill_2
XFILLER_22_964 VPWR VGND sg13g2_decap_8
X_5878_ VPWR _0168_ _1497_ VGND sg13g2_inv_1
X_4829_ net1134 net1066 _0552_ VPWR VGND sg13g2_nor2b_1
XFILLER_4_128 VPWR VGND sg13g2_fill_1
XFILLER_1_802 VPWR VGND sg13g2_decap_8
XFILLER_0_301 VPWR VGND sg13g2_decap_8
XFILLER_1_879 VPWR VGND sg13g2_decap_8
XFILLER_49_828 VPWR VGND sg13g2_decap_8
XFILLER_17_714 VPWR VGND sg13g2_decap_4
XFILLER_1_1028 VPWR VGND sg13g2_fill_1
XFILLER_16_202 VPWR VGND sg13g2_fill_2
XFILLER_29_596 VPWR VGND sg13g2_decap_8
XFILLER_17_94 VPWR VGND sg13g2_fill_2
XFILLER_13_942 VPWR VGND sg13g2_decap_8
XFILLER_31_238 VPWR VGND sg13g2_decap_4
X_6203__53 VPWR VGND net53 sg13g2_tiehi
XFILLER_9_957 VPWR VGND sg13g2_decap_8
XFILLER_4_673 VPWR VGND sg13g2_fill_1
XFILLER_3_161 VPWR VGND sg13g2_decap_8
X_3160_ net1001 net1066 _1611_ VPWR VGND sg13g2_nor2b_1
Xhold1 s0.genblk1\[1\].modules.bubble VPWR VGND net297 sg13g2_dlygate4sd3_1
XFILLER_48_850 VPWR VGND sg13g2_decap_8
XFILLER_35_588 VPWR VGND sg13g2_decap_8
X_5801_ VGND VPWR _1366_ _1421_ _1427_ net1279 sg13g2_a21oi_1
X_6162__111 VPWR VGND net111 sg13g2_tiehi
XFILLER_16_780 VPWR VGND sg13g2_decap_4
X_5732_ s0.data_out\[8\]\[1\] s0.data_out\[9\]\[1\] net1041 _1365_ VPWR VGND sg13g2_mux2_1
X_3993_ net1261 _2365_ _2366_ VPWR VGND sg13g2_and2_1
XFILLER_31_772 VPWR VGND sg13g2_decap_4
X_5663_ s0.data_out\[10\]\[3\] s0.data_out\[9\]\[3\] net1041 _1308_ VPWR VGND sg13g2_mux2_1
X_4614_ VGND VPWR net1157 net341 _0356_ _0355_ sg13g2_a21oi_1
X_5594_ s0.data_out\[9\]\[1\] s0.data_out\[10\]\[1\] net1084 _1246_ VPWR VGND sg13g2_mux2_1
X_4545_ _0294_ _0295_ _0296_ VPWR VGND sg13g2_nor2_1
X_4476_ net1287 VPWR _2794_ VGND net927 _2793_ sg13g2_o21ai_1
Xfanout914 _2471_ net914 VPWR VGND sg13g2_buf_8
Xfanout925 _2461_ net925 VPWR VGND sg13g2_buf_8
X_3427_ _1849_ _1852_ net1311 _1853_ VPWR VGND sg13g2_nand3_1
X_6215_ net149 VGND VPWR _0265_ s0.data_out\[0\]\[3\] clknet_leaf_7_clk sg13g2_dfrbpq_1
Xfanout958 s0.valid_out\[1\][0] net958 VPWR VGND sg13g2_buf_8
X_6146_ net128 VGND VPWR _0196_ s0.data_out\[6\]\[6\] clknet_leaf_12_clk sg13g2_dfrbpq_2
X_3358_ _1791_ net998 net538 VPWR VGND sg13g2_nand2_1
Xfanout947 net948 net947 VPWR VGND sg13g2_buf_8
Xfanout936 _2453_ net936 VPWR VGND sg13g2_buf_1
Xfanout969 net970 net969 VPWR VGND sg13g2_buf_2
X_6077_ net202 VGND VPWR _0127_ s0.data_out\[11\]\[4\] clknet_leaf_21_clk sg13g2_dfrbpq_2
X_3289_ net991 net1066 _1728_ VPWR VGND sg13g2_nor2b_1
X_5028_ _0733_ net1132 net598 VPWR VGND sg13g2_nand2_1
XFILLER_13_249 VPWR VGND sg13g2_decap_4
XFILLER_10_901 VPWR VGND sg13g2_fill_2
XFILLER_16_1014 VPWR VGND sg13g2_decap_8
XFILLER_6_905 VPWR VGND sg13g2_decap_8
XFILLER_5_426 VPWR VGND sg13g2_decap_8
XFILLER_10_989 VPWR VGND sg13g2_decap_8
X_6139__135 VPWR VGND net135 sg13g2_tiehi
XFILLER_49_625 VPWR VGND sg13g2_decap_8
XFILLER_1_676 VPWR VGND sg13g2_decap_8
XFILLER_17_500 VPWR VGND sg13g2_fill_1
XFILLER_28_93 VPWR VGND sg13g2_fill_1
XFILLER_44_341 VPWR VGND sg13g2_decap_8
XFILLER_44_330 VPWR VGND sg13g2_fill_2
X_6146__128 VPWR VGND net128 sg13g2_tiehi
XFILLER_45_886 VPWR VGND sg13g2_decap_8
XFILLER_17_599 VPWR VGND sg13g2_fill_1
XFILLER_20_709 VPWR VGND sg13g2_decap_8
XFILLER_8_220 VPWR VGND sg13g2_fill_2
XFILLER_5_993 VPWR VGND sg13g2_decap_8
X_4330_ _2662_ net931 _2661_ VPWR VGND sg13g2_nand2_1
X_4261_ VGND VPWR _2601_ _2598_ net1239 sg13g2_or2_1
X_6000_ net285 VGND VPWR _0050_ s0.valid_out\[17\][0] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3212_ _1657_ net1012 _1656_ VPWR VGND sg13g2_nand2b_1
X_4192_ net1202 VPWR _2537_ VGND _2535_ _2536_ sg13g2_o21ai_1
XFILLER_39_146 VPWR VGND sg13g2_fill_2
X_3143_ net1001 s0.data_out\[6\]\[0\] _1596_ VPWR VGND sg13g2_and2_1
XFILLER_39_1014 VPWR VGND sg13g2_decap_8
X_3976_ VGND VPWR net942 _2348_ _2349_ _2308_ sg13g2_a21oi_1
X_5715_ VPWR _1351_ _1350_ VGND sg13g2_inv_1
XFILLER_10_219 VPWR VGND sg13g2_decap_4
X_5646_ net1347 VPWR _1292_ VGND net934 _1291_ sg13g2_o21ai_1
XFILLER_40_39 VPWR VGND sg13g2_fill_1
Xhold220 _2116_ VPWR VGND net516 sg13g2_dlygate4sd3_1
XFILLER_3_908 VPWR VGND sg13g2_decap_8
X_5577_ VPWR _1232_ _1231_ VGND sg13g2_inv_1
Xhold242 s0.data_out\[5\]\[6\] VPWR VGND net538 sg13g2_dlygate4sd3_1
XFILLER_2_407 VPWR VGND sg13g2_decap_8
X_4528_ _0281_ net1183 _0280_ VPWR VGND sg13g2_nand2b_1
Xhold253 _0812_ VPWR VGND net549 sg13g2_dlygate4sd3_1
Xhold231 s0.data_out\[11\]\[6\] VPWR VGND net527 sg13g2_dlygate4sd3_1
Xhold264 s0.data_out\[20\]\[3\] VPWR VGND net560 sg13g2_dlygate4sd3_1
Xhold286 s0.data_out\[17\]\[5\] VPWR VGND net582 sg13g2_dlygate4sd3_1
X_4459_ net1170 net1057 _2779_ VPWR VGND sg13g2_nor2b_1
Xhold275 _0345_ VPWR VGND net571 sg13g2_dlygate4sd3_1
XFILLER_49_59 VPWR VGND sg13g2_fill_2
Xhold297 s0.data_new_delayed\[7\] VPWR VGND net593 sg13g2_dlygate4sd3_1
X_6129_ net146 VGND VPWR _0179_ s0.data_out\[7\]\[1\] clknet_leaf_23_clk sg13g2_dfrbpq_2
XFILLER_45_138 VPWR VGND sg13g2_fill_1
XFILLER_42_812 VPWR VGND sg13g2_fill_1
XFILLER_14_40 VPWR VGND sg13g2_fill_2
XFILLER_10_753 VPWR VGND sg13g2_fill_2
XFILLER_2_952 VPWR VGND sg13g2_decap_8
X_6152__121 VPWR VGND net121 sg13g2_tiehi
XFILLER_49_422 VPWR VGND sg13g2_decap_8
XFILLER_49_499 VPWR VGND sg13g2_decap_8
XFILLER_17_341 VPWR VGND sg13g2_fill_2
XFILLER_44_193 VPWR VGND sg13g2_decap_8
X_3830_ VPWR _0243_ _2217_ VGND sg13g2_inv_1
XFILLER_20_506 VPWR VGND sg13g2_fill_2
XFILLER_33_867 VPWR VGND sg13g2_fill_1
X_3761_ _2156_ _2157_ _2158_ VPWR VGND sg13g2_nor2_1
X_5500_ _1160_ net481 net1097 VPWR VGND sg13g2_nand2b_1
XFILLER_9_584 VPWR VGND sg13g2_fill_2
X_3692_ net971 VPWR _2093_ VGND _2091_ _2092_ sg13g2_o21ai_1
X_5431_ _1100_ net1098 net541 VPWR VGND sg13g2_nand2_1
X_5362_ VGND VPWR _0978_ _1034_ _1035_ net1103 sg13g2_a21oi_1
X_4313_ _2647_ net475 net1199 VPWR VGND sg13g2_nand2b_1
X_5293_ VGND VPWR _0974_ _0972_ net1242 sg13g2_or2_1
X_4244_ _2584_ net1198 net560 VPWR VGND sg13g2_nand2_1
XFILLER_19_29 VPWR VGND sg13g2_decap_8
X_4175_ net1190 net1069 _2522_ VPWR VGND sg13g2_nor2b_1
X_3126_ VGND VPWR _1583_ net1209 net307 sg13g2_or2_1
XFILLER_28_617 VPWR VGND sg13g2_fill_2
XFILLER_42_108 VPWR VGND sg13g2_fill_2
XFILLER_24_812 VPWR VGND sg13g2_decap_8
XFILLER_35_171 VPWR VGND sg13g2_fill_2
X_3959_ VGND VPWR _2256_ _2333_ _2334_ net952 sg13g2_a21oi_1
XFILLER_13_1028 VPWR VGND sg13g2_fill_1
X_5629_ net1038 net1055 _1277_ VPWR VGND sg13g2_nor2b_1
X_6190__80 VPWR VGND net80 sg13g2_tiehi
XFILLER_47_948 VPWR VGND sg13g2_decap_8
XFILLER_46_414 VPWR VGND sg13g2_fill_1
XFILLER_27_650 VPWR VGND sg13g2_decap_8
XFILLER_14_333 VPWR VGND sg13g2_decap_4
XFILLER_14_399 VPWR VGND sg13g2_decap_8
XFILLER_30_815 VPWR VGND sg13g2_decap_4
XFILLER_30_859 VPWR VGND sg13g2_fill_2
XFILLER_6_554 VPWR VGND sg13g2_decap_4
XFILLER_6_521 VPWR VGND sg13g2_decap_8
XFILLER_10_594 VPWR VGND sg13g2_fill_1
XFILLER_44_7 VPWR VGND sg13g2_fill_1
XFILLER_29_1002 VPWR VGND sg13g2_decap_8
XFILLER_49_241 VPWR VGND sg13g2_decap_8
XFILLER_49_252 VPWR VGND sg13g2_decap_8
XFILLER_38_926 VPWR VGND sg13g2_decap_8
XFILLER_37_414 VPWR VGND sg13g2_decap_4
X_5980_ net35 VGND VPWR _0030_ s0.data_out\[19\]\[3\] clknet_leaf_37_clk sg13g2_dfrbpq_2
XFILLER_46_992 VPWR VGND sg13g2_decap_8
X_4931_ VGND VPWR _0646_ net1130 net378 sg13g2_or2_1
X_4862_ net1317 VPWR _0581_ VGND net923 _0580_ sg13g2_o21ai_1
X_3813_ _2202_ VPWR _2203_ VGND net1297 net446 sg13g2_o21ai_1
X_4793_ _0522_ _0505_ _0504_ VPWR VGND sg13g2_nand2b_1
X_3744_ s0.data_out\[3\]\[6\] s0.data_out\[2\]\[6\] net967 _2141_ VPWR VGND sg13g2_mux2_1
X_3675_ net959 net1068 _2078_ VPWR VGND sg13g2_nor2b_1
X_5414_ _1083_ net1097 net540 VPWR VGND sg13g2_nand2_1
XFILLER_0_719 VPWR VGND sg13g2_decap_8
X_5345_ _1020_ s0.data_out\[11\]\[2\] net1109 VPWR VGND sg13g2_nand2b_1
X_5276_ VGND VPWR _0896_ _0951_ _0957_ net1279 sg13g2_a21oi_1
X_4227_ net1203 _2566_ _2567_ _2568_ VPWR VGND sg13g2_nor3_1
X_4158_ s0.was_valid_out\[20\][0] net1200 _2508_ VPWR VGND sg13g2_nor2_1
X_3109_ VGND VPWR net1016 _1565_ _1566_ _1508_ sg13g2_a21oi_1
X_4089_ VPWR _2448_ net1093 VGND sg13g2_inv_1
XFILLER_37_992 VPWR VGND sg13g2_decap_8
XFILLER_12_859 VPWR VGND sg13g2_decap_4
XFILLER_20_870 VPWR VGND sg13g2_fill_2
X_6003__282 VPWR VGND net282 sg13g2_tiehi
XFILLER_3_568 VPWR VGND sg13g2_fill_2
XFILLER_3_557 VPWR VGND sg13g2_decap_8
Xfanout1314 net1315 net1314 VPWR VGND sg13g2_buf_1
Xfanout1303 net1316 net1303 VPWR VGND sg13g2_buf_8
Xfanout1325 net1326 net1325 VPWR VGND sg13g2_buf_8
Xfanout1336 net1337 net1336 VPWR VGND sg13g2_buf_8
Xfanout1347 net1348 net1347 VPWR VGND sg13g2_buf_2
XFILLER_47_745 VPWR VGND sg13g2_decap_8
XFILLER_4_1026 VPWR VGND sg13g2_fill_2
X_5969__47 VPWR VGND net47 sg13g2_tiehi
XFILLER_43_940 VPWR VGND sg13g2_decap_8
XFILLER_36_93 VPWR VGND sg13g2_fill_2
X_6010__275 VPWR VGND net275 sg13g2_tiehi
XFILLER_14_185 VPWR VGND sg13g2_fill_1
XFILLER_7_852 VPWR VGND sg13g2_fill_1
XFILLER_10_391 VPWR VGND sg13g2_decap_8
X_3460_ _1881_ VPWR _1882_ VGND _1877_ _1880_ sg13g2_o21ai_1
X_3391_ VGND VPWR _1822_ net989 net353 sg13g2_or2_1
X_5130_ net1333 VPWR _0824_ VGND net937 _0823_ sg13g2_o21ai_1
X_5061_ VPWR _0764_ _0763_ VGND sg13g2_inv_1
X_4012_ VGND VPWR net943 _2384_ _2385_ _2329_ sg13g2_a21oi_1
XFILLER_38_778 VPWR VGND sg13g2_decap_4
XFILLER_37_244 VPWR VGND sg13g2_fill_1
XFILLER_25_406 VPWR VGND sg13g2_fill_1
X_5963_ net54 VGND VPWR _0013_ s0.was_valid_out\[20\][0] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_4914_ _0564_ _0629_ net1258 _0631_ VPWR VGND sg13g2_nand3_1
X_5894_ VPWR _0170_ _1511_ VGND sg13g2_inv_1
XFILLER_34_984 VPWR VGND sg13g2_decap_8
X_4845_ net1136 net1059 _0566_ VPWR VGND sg13g2_nor2b_1
X_4776_ VGND VPWR _0505_ _0503_ net1233 sg13g2_or2_1
XFILLER_21_667 VPWR VGND sg13g2_decap_4
XFILLER_21_689 VPWR VGND sg13g2_fill_1
X_3727_ _2069_ _2123_ net1275 _2124_ VPWR VGND sg13g2_nand3_1
X_3658_ net959 s0.data_out\[2\]\[0\] _2063_ VPWR VGND sg13g2_and2_1
X_3589_ _1998_ VPWR _1999_ VGND _1994_ _1997_ sg13g2_o21ai_1
XFILLER_0_516 VPWR VGND sg13g2_decap_8
X_5328_ net1220 _1000_ _0110_ VPWR VGND sg13g2_nor2_1
X_5259_ net1338 VPWR _0941_ VGND net936 _0940_ sg13g2_o21ai_1
XFILLER_29_712 VPWR VGND sg13g2_decap_8
XFILLER_44_715 VPWR VGND sg13g2_decap_8
XFILLER_17_907 VPWR VGND sg13g2_fill_1
XFILLER_43_225 VPWR VGND sg13g2_fill_1
XFILLER_44_759 VPWR VGND sg13g2_fill_1
XFILLER_19_1001 VPWR VGND sg13g2_decap_8
XFILLER_43_269 VPWR VGND sg13g2_fill_1
XFILLER_24_450 VPWR VGND sg13g2_fill_2
XFILLER_11_100 VPWR VGND sg13g2_fill_1
XFILLER_40_987 VPWR VGND sg13g2_decap_8
XFILLER_12_678 VPWR VGND sg13g2_fill_1
XFILLER_12_689 VPWR VGND sg13g2_fill_2
XFILLER_4_844 VPWR VGND sg13g2_decap_8
XFILLER_3_387 VPWR VGND sg13g2_decap_4
XFILLER_0_0 VPWR VGND sg13g2_decap_8
Xfanout1122 net1123 net1122 VPWR VGND sg13g2_buf_2
Xfanout1100 net1104 net1100 VPWR VGND sg13g2_buf_8
Xfanout1111 s0.valid_out\[12\][0] net1111 VPWR VGND sg13g2_buf_8
Xfanout1155 net1157 net1155 VPWR VGND sg13g2_buf_8
Xfanout1144 net1145 net1144 VPWR VGND sg13g2_buf_2
Xfanout1133 s0.valid_out\[14\][0] net1133 VPWR VGND sg13g2_buf_8
XFILLER_47_520 VPWR VGND sg13g2_decap_8
Xfanout1199 net1201 net1199 VPWR VGND sg13g2_buf_1
Xfanout1177 s0.valid_out\[18\][0] net1177 VPWR VGND sg13g2_buf_8
Xfanout1188 net1189 net1188 VPWR VGND sg13g2_buf_8
Xfanout1166 s0.valid_out\[17\][0] net1166 VPWR VGND sg13g2_buf_8
XFILLER_35_715 VPWR VGND sg13g2_decap_4
XFILLER_35_737 VPWR VGND sg13g2_decap_8
XFILLER_15_450 VPWR VGND sg13g2_fill_2
XFILLER_15_461 VPWR VGND sg13g2_fill_1
X_4630_ _0371_ net1169 _0370_ VPWR VGND sg13g2_nand2b_1
XFILLER_30_442 VPWR VGND sg13g2_fill_1
XFILLER_8_75 VPWR VGND sg13g2_decap_4
XFILLER_8_53 VPWR VGND sg13g2_fill_2
XFILLER_30_475 VPWR VGND sg13g2_fill_1
X_4561_ _0309_ VPWR _0310_ VGND net1301 net460 sg13g2_o21ai_1
X_3512_ VGND VPWR _1933_ net1208 net318 sg13g2_or2_1
X_4492_ _2808_ net1174 net493 VPWR VGND sg13g2_nand2_1
X_3443_ _1863_ _1866_ net1314 _1867_ VPWR VGND sg13g2_nand3_1
X_6162_ net111 VGND VPWR _0212_ s0.was_valid_out\[4\][0] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_5113_ VGND VPWR net1114 s0.data_out\[13\]\[5\] _0809_ _0808_ sg13g2_a21oi_1
XFILLER_33_0 VPWR VGND sg13g2_decap_4
X_3374_ _1806_ _1741_ net1258 _1807_ VPWR VGND sg13g2_a21o_1
X_6093_ net185 VGND VPWR _0143_ s0.shift_out\[10\][0] clknet_leaf_19_clk sg13g2_dfrbpq_2
X_5044_ VGND VPWR net1125 _0748_ _0749_ _0689_ sg13g2_a21oi_1
XFILLER_38_586 VPWR VGND sg13g2_fill_2
XFILLER_41_718 VPWR VGND sg13g2_decap_8
X_5946_ _1560_ _1559_ net1243 _1555_ net1237 VPWR VGND sg13g2_a22oi_1
X_5956__61 VPWR VGND net61 sg13g2_tiehi
X_5877_ _1496_ VPWR _1497_ VGND _1492_ _1495_ sg13g2_o21ai_1
XFILLER_33_280 VPWR VGND sg13g2_decap_8
X_4828_ net1134 s0.data_out\[15\]\[2\] _0551_ VPWR VGND sg13g2_and2_1
X_4759_ _0480_ VPWR _0488_ VGND net1277 _0483_ sg13g2_o21ai_1
XFILLER_49_807 VPWR VGND sg13g2_decap_8
XFILLER_1_858 VPWR VGND sg13g2_decap_8
X_6000__285 VPWR VGND net285 sg13g2_tiehi
XFILLER_0_379 VPWR VGND sg13g2_decap_8
XFILLER_12_420 VPWR VGND sg13g2_decap_4
XFILLER_31_228 VPWR VGND sg13g2_fill_1
XFILLER_9_936 VPWR VGND sg13g2_decap_8
XFILLER_12_442 VPWR VGND sg13g2_decap_4
XFILLER_13_998 VPWR VGND sg13g2_decap_8
Xhold2 s0.genblk1\[13\].modules.bubble VPWR VGND net298 sg13g2_dlygate4sd3_1
XFILLER_0_880 VPWR VGND sg13g2_decap_8
XFILLER_35_501 VPWR VGND sg13g2_fill_2
X_5800_ net1283 _1425_ _1426_ VPWR VGND sg13g2_nor2b_1
X_3992_ VGND VPWR net951 _2364_ _2365_ _2313_ sg13g2_a21oi_1
X_5731_ VPWR _0154_ _1364_ VGND sg13g2_inv_1
XFILLER_15_291 VPWR VGND sg13g2_fill_2
X_5662_ _1298_ VPWR _1307_ VGND net1278 _1302_ sg13g2_o21ai_1
X_5953__64 VPWR VGND net64 sg13g2_tiehi
X_4613_ net1157 net1046 _0355_ VPWR VGND sg13g2_nor2b_1
X_5593_ VPWR _0135_ _1245_ VGND sg13g2_inv_1
X_4544_ net1226 net1163 _0295_ VPWR VGND sg13g2_nor2b_1
XFILLER_7_490 VPWR VGND sg13g2_fill_2
X_4475_ VGND VPWR net1170 s0.data_out\[18\]\[6\] _2793_ _2792_ sg13g2_a21oi_1
X_6214_ net162 VGND VPWR _0264_ s0.data_out\[0\]\[2\] clknet_leaf_7_clk sg13g2_dfrbpq_1
Xfanout915 _2470_ net915 VPWR VGND sg13g2_buf_8
X_3426_ net990 VPWR _1852_ VGND _1850_ _1851_ sg13g2_o21ai_1
X_6145_ net129 VGND VPWR _0195_ s0.data_out\[6\]\[5\] clknet_leaf_17_clk sg13g2_dfrbpq_2
Xfanout948 s0.valid_out\[0\][0] net948 VPWR VGND sg13g2_buf_8
X_3357_ VGND VPWR net1007 _1789_ _1790_ _1762_ sg13g2_a21oi_1
Xfanout926 _2460_ net926 VPWR VGND sg13g2_buf_8
Xfanout937 _2452_ net937 VPWR VGND sg13g2_buf_8
X_6076_ net203 VGND VPWR _0126_ s0.data_out\[11\]\[3\] clknet_leaf_25_clk sg13g2_dfrbpq_2
Xfanout959 net960 net959 VPWR VGND sg13g2_buf_8
X_5027_ VGND VPWR net1139 _0731_ _0732_ _0701_ sg13g2_a21oi_1
X_3288_ VGND VPWR _1650_ _1726_ _1727_ net1000 sg13g2_a21oi_1
XFILLER_26_534 VPWR VGND sg13g2_fill_2
XFILLER_14_729 VPWR VGND sg13g2_fill_1
X_5929_ VPWR VGND _1478_ net1283 _1542_ net1278 _1543_ _1539_ sg13g2_a221oi_1
XFILLER_10_968 VPWR VGND sg13g2_decap_8
XFILLER_49_604 VPWR VGND sg13g2_decap_8
XFILLER_1_655 VPWR VGND sg13g2_decap_8
XFILLER_0_165 VPWR VGND sg13g2_decap_8
XFILLER_45_865 VPWR VGND sg13g2_decap_8
XFILLER_32_515 VPWR VGND sg13g2_fill_2
XFILLER_13_740 VPWR VGND sg13g2_fill_2
XFILLER_12_250 VPWR VGND sg13g2_decap_4
XFILLER_9_766 VPWR VGND sg13g2_decap_8
X_6081__198 VPWR VGND net198 sg13g2_tiehi
XFILLER_8_265 VPWR VGND sg13g2_decap_4
XFILLER_5_972 VPWR VGND sg13g2_decap_8
XFILLER_5_54 VPWR VGND sg13g2_fill_1
X_4260_ net1231 _2594_ _2600_ VPWR VGND sg13g2_nor2_1
X_4191_ net1190 net1061 _2536_ VPWR VGND sg13g2_nor2b_1
X_3211_ VGND VPWR net1001 _1655_ _1656_ _1604_ sg13g2_a21oi_1
X_3142_ _1595_ net917 _1594_ VPWR VGND sg13g2_nand2_1
XFILLER_23_537 VPWR VGND sg13g2_fill_2
XFILLER_23_559 VPWR VGND sg13g2_fill_2
X_3975_ _2347_ VPWR _2348_ VGND net946 _2493_ sg13g2_o21ai_1
X_5714_ _1348_ _1349_ _1350_ VPWR VGND sg13g2_nor2_1
X_5645_ VGND VPWR net1038 s0.data_out\[9\]\[7\] _1291_ _1290_ sg13g2_a21oi_1
Xhold210 s0.data_out\[10\]\[2\] VPWR VGND net506 sg13g2_dlygate4sd3_1
X_5576_ _1229_ _1230_ _1231_ VPWR VGND sg13g2_nor2_1
Xhold243 s0.data_out\[6\]\[5\] VPWR VGND net539 sg13g2_dlygate4sd3_1
Xhold221 s0.data_out\[7\]\[7\] VPWR VGND net517 sg13g2_dlygate4sd3_1
Xhold232 s0.data_out\[12\]\[1\] VPWR VGND net528 sg13g2_dlygate4sd3_1
X_4527_ VGND VPWR net1170 _0279_ _0280_ _2779_ sg13g2_a21oi_1
Xhold254 s0.data_out\[16\]\[3\] VPWR VGND net550 sg13g2_dlygate4sd3_1
Xhold265 _2660_ VPWR VGND net561 sg13g2_dlygate4sd3_1
Xhold276 s0.data_out\[17\]\[6\] VPWR VGND net572 sg13g2_dlygate4sd3_1
X_4458_ net1170 s0.data_out\[18\]\[4\] _2778_ VPWR VGND sg13g2_and2_1
Xhold287 _0462_ VPWR VGND net583 sg13g2_dlygate4sd3_1
XFILLER_49_49 VPWR VGND sg13g2_fill_2
Xhold298 s0.data_out\[12\]\[7\] VPWR VGND net594 sg13g2_dlygate4sd3_1
X_3409_ net981 net1070 _1837_ VPWR VGND sg13g2_nor2b_1
X_4389_ _2717_ _2716_ net1239 _2712_ net1231 VPWR VGND sg13g2_a22oi_1
X_6128_ net147 VGND VPWR _0178_ s0.data_out\[7\]\[0\] clknet_leaf_23_clk sg13g2_dfrbpq_2
X_6059_ net222 VGND VPWR net409 s0.was_valid_out\[12\][0] clknet_leaf_26_clk sg13g2_dfrbpq_2
XFILLER_27_865 VPWR VGND sg13g2_decap_4
XFILLER_14_515 VPWR VGND sg13g2_decap_8
XFILLER_41_345 VPWR VGND sg13g2_decap_8
XFILLER_10_732 VPWR VGND sg13g2_fill_1
XFILLER_6_725 VPWR VGND sg13g2_fill_2
XFILLER_5_213 VPWR VGND sg13g2_fill_2
XFILLER_30_51 VPWR VGND sg13g2_fill_2
XFILLER_2_931 VPWR VGND sg13g2_decap_8
XFILLER_49_401 VPWR VGND sg13g2_decap_8
XFILLER_7_1013 VPWR VGND sg13g2_decap_8
XFILLER_49_478 VPWR VGND sg13g2_decap_8
XFILLER_36_106 VPWR VGND sg13g2_fill_1
XFILLER_32_345 VPWR VGND sg13g2_decap_4
XFILLER_20_529 VPWR VGND sg13g2_fill_1
X_3760_ net1262 _2133_ _2157_ VPWR VGND sg13g2_nor2_1
XFILLER_9_596 VPWR VGND sg13g2_fill_2
X_5430_ _1099_ net1256 _1098_ VPWR VGND sg13g2_nand2_1
X_3691_ net960 net1058 _2092_ VPWR VGND sg13g2_nor2b_1
X_5361_ _1034_ net330 net1110 VPWR VGND sg13g2_nand2b_1
XFILLER_5_780 VPWR VGND sg13g2_fill_2
X_4312_ VPWR _0016_ _2646_ VGND sg13g2_inv_1
X_5292_ _0973_ _0972_ net1242 _0968_ net1236 VPWR VGND sg13g2_a22oi_1
X_4243_ VPWR VGND _2581_ _2582_ _2577_ net1211 _2583_ _2573_ sg13g2_a221oi_1
X_4174_ net1190 s0.data_out\[20\]\[1\] _2521_ VPWR VGND sg13g2_and2_1
X_3125_ _1471_ _1580_ _1581_ _1582_ VPWR VGND sg13g2_nor3_1
X_6129__146 VPWR VGND net146 sg13g2_tiehi
XFILLER_24_835 VPWR VGND sg13g2_decap_8
X_3958_ _2333_ net351 net956 VPWR VGND sg13g2_nand2b_1
X_3889_ VGND VPWR _2212_ _2271_ _2274_ net1247 sg13g2_a21oi_1
X_5628_ net919 _2490_ _1276_ VPWR VGND sg13g2_nor2_1
X_5559_ _1215_ net1080 _1162_ _1216_ VPWR VGND sg13g2_a21o_1
X_6136__139 VPWR VGND net139 sg13g2_tiehi
XFILLER_47_927 VPWR VGND sg13g2_decap_8
XFILLER_19_629 VPWR VGND sg13g2_decap_4
XFILLER_14_312 VPWR VGND sg13g2_fill_1
XFILLER_15_868 VPWR VGND sg13g2_decap_8
XFILLER_41_50 VPWR VGND sg13g2_decap_4
XFILLER_10_540 VPWR VGND sg13g2_fill_2
XFILLER_49_275 VPWR VGND sg13g2_decap_8
XFILLER_49_297 VPWR VGND sg13g2_decap_8
XFILLER_2_88 VPWR VGND sg13g2_decap_4
XFILLER_2_99 VPWR VGND sg13g2_fill_1
XFILLER_46_971 VPWR VGND sg13g2_decap_8
XFILLER_18_662 VPWR VGND sg13g2_fill_2
XFILLER_45_481 VPWR VGND sg13g2_fill_2
X_4930_ VGND VPWR _0645_ _0644_ _0643_ sg13g2_or2_1
XFILLER_17_161 VPWR VGND sg13g2_decap_4
X_4861_ VGND VPWR net1136 s0.data_out\[15\]\[6\] _0580_ _0579_ sg13g2_a21oi_1
XFILLER_21_816 VPWR VGND sg13g2_decap_8
XFILLER_32_164 VPWR VGND sg13g2_decap_8
X_3812_ _2198_ _2201_ net1297 _2202_ VPWR VGND sg13g2_nand3_1
X_4792_ _0521_ _0515_ _0520_ VPWR VGND sg13g2_nand2_1
X_3743_ _2140_ net966 net491 VPWR VGND sg13g2_nand2_1
XFILLER_20_359 VPWR VGND sg13g2_fill_1
X_3674_ net959 net611 _2077_ VPWR VGND sg13g2_and2_1
X_5413_ VPWR VGND net1265 _1076_ _1081_ net1270 _1082_ _1065_ sg13g2_a221oi_1
X_5344_ VPWR _0112_ net529 VGND sg13g2_inv_1
X_5275_ net1282 _0955_ _0956_ VPWR VGND sg13g2_nor2b_1
X_4226_ net1207 s0.data_out\[20\]\[7\] _2567_ VPWR VGND sg13g2_nor2_1
XFILLER_29_905 VPWR VGND sg13g2_fill_1
X_4157_ _2505_ VPWR _2507_ VGND net1205 _2506_ sg13g2_o21ai_1
X_3108_ s0.data_out\[8\]\[4\] s0.data_out\[7\]\[4\] net1021 _1565_ VPWR VGND sg13g2_mux2_1
XFILLER_37_971 VPWR VGND sg13g2_decap_8
X_5978__37 VPWR VGND net37 sg13g2_tiehi
X_4088_ VPWR _2447_ net323 VGND sg13g2_inv_1
XFILLER_28_459 VPWR VGND sg13g2_fill_1
XFILLER_24_643 VPWR VGND sg13g2_decap_4
XFILLER_24_676 VPWR VGND sg13g2_decap_8
X_6142__132 VPWR VGND net132 sg13g2_tiehi
XFILLER_20_860 VPWR VGND sg13g2_fill_1
Xfanout1304 net1305 net1304 VPWR VGND sg13g2_buf_8
Xfanout1337 net1339 net1337 VPWR VGND sg13g2_buf_8
Xfanout1315 net1316 net1315 VPWR VGND sg13g2_buf_8
Xfanout1326 net1349 net1326 VPWR VGND sg13g2_buf_8
Xfanout1348 net1349 net1348 VPWR VGND sg13g2_buf_8
XFILLER_4_1005 VPWR VGND sg13g2_decap_8
XFILLER_47_724 VPWR VGND sg13g2_decap_8
XFILLER_15_610 VPWR VGND sg13g2_decap_8
XFILLER_28_993 VPWR VGND sg13g2_decap_8
XFILLER_43_996 VPWR VGND sg13g2_decap_8
XFILLER_6_341 VPWR VGND sg13g2_decap_8
X_3390_ VGND VPWR _1821_ _1820_ _1819_ sg13g2_or2_1
X_5060_ VGND VPWR _2449_ net1119 _0763_ _0762_ sg13g2_a21oi_1
X_4011_ s0.data_out\[1\]\[5\] s0.data_out\[0\]\[5\] net947 _2384_ VPWR VGND sg13g2_mux2_1
XFILLER_38_713 VPWR VGND sg13g2_fill_2
XFILLER_38_746 VPWR VGND sg13g2_fill_2
XFILLER_37_267 VPWR VGND sg13g2_fill_2
X_5962_ net55 VGND VPWR _0012_ s0.genblk1\[20\].modules.bubble clknet_leaf_2_clk sg13g2_dfrbpq_1
X_4913_ VGND VPWR _0564_ _0629_ _0630_ net1258 sg13g2_a21oi_1
XFILLER_34_963 VPWR VGND sg13g2_decap_8
X_5893_ _1510_ VPWR _1511_ VGND net1330 net350 sg13g2_o21ai_1
X_4844_ net1137 s0.data_out\[15\]\[4\] _0565_ VPWR VGND sg13g2_and2_1
XFILLER_20_101 VPWR VGND sg13g2_fill_2
XFILLER_32_19 VPWR VGND sg13g2_fill_2
X_4775_ _0504_ _0503_ net1233 _0499_ net1240 VPWR VGND sg13g2_a22oi_1
XFILLER_20_189 VPWR VGND sg13g2_decap_4
X_3726_ _2123_ net971 _2122_ VPWR VGND sg13g2_nand2b_1
X_3657_ _2062_ net932 _2061_ VPWR VGND sg13g2_nand2_1
X_3588_ VGND VPWR _1998_ net535 net1313 sg13g2_or2_1
X_5327_ _1004_ _1005_ _0109_ VPWR VGND sg13g2_nor2_1
X_5258_ VGND VPWR net1107 s0.data_out\[12\]\[7\] _0940_ _0939_ sg13g2_a21oi_1
X_5189_ _0878_ _0879_ _0880_ VPWR VGND sg13g2_nor2_1
X_4209_ net361 s0.valid_out\[21\][0] _2552_ VPWR VGND sg13g2_nor2b_1
XFILLER_25_930 VPWR VGND sg13g2_fill_2
XFILLER_25_985 VPWR VGND sg13g2_decap_8
XFILLER_12_624 VPWR VGND sg13g2_fill_1
XFILLER_40_966 VPWR VGND sg13g2_decap_8
XFILLER_7_116 VPWR VGND sg13g2_fill_1
XFILLER_20_690 VPWR VGND sg13g2_decap_8
XFILLER_4_823 VPWR VGND sg13g2_decap_8
Xfanout1112 net1113 net1112 VPWR VGND sg13g2_buf_2
Xfanout1101 net1104 net1101 VPWR VGND sg13g2_buf_1
Xfanout1156 net1157 net1156 VPWR VGND sg13g2_buf_1
Xfanout1134 net1135 net1134 VPWR VGND sg13g2_buf_8
Xfanout1145 net1147 net1145 VPWR VGND sg13g2_buf_1
Xfanout1123 net1124 net1123 VPWR VGND sg13g2_buf_1
Xfanout1167 net1168 net1167 VPWR VGND sg13g2_buf_2
Xfanout1178 net1179 net1178 VPWR VGND sg13g2_buf_2
Xfanout1189 net337 net1189 VPWR VGND sg13g2_buf_8
XFILLER_19_201 VPWR VGND sg13g2_fill_2
XFILLER_19_212 VPWR VGND sg13g2_fill_2
XFILLER_47_565 VPWR VGND sg13g2_fill_2
XFILLER_19_245 VPWR VGND sg13g2_decap_8
XFILLER_16_941 VPWR VGND sg13g2_fill_1
XFILLER_16_952 VPWR VGND sg13g2_fill_2
XFILLER_15_440 VPWR VGND sg13g2_fill_2
X_5965__51 VPWR VGND net51 sg13g2_tiehi
XFILLER_30_410 VPWR VGND sg13g2_fill_1
X_4560_ _0305_ _0308_ net1301 _0309_ VPWR VGND sg13g2_nand3_1
XFILLER_31_999 VPWR VGND sg13g2_decap_8
XFILLER_11_690 VPWR VGND sg13g2_fill_1
X_3511_ _1821_ _1930_ _1931_ _1932_ VPWR VGND sg13g2_nor3_1
XFILLER_7_672 VPWR VGND sg13g2_decap_8
X_4491_ _2763_ VPWR _2807_ VGND net926 _2806_ sg13g2_o21ai_1
X_3442_ net994 VPWR _1866_ VGND _1864_ _1865_ sg13g2_o21ai_1
X_6161_ net112 VGND VPWR _0211_ s0.genblk1\[4\].modules.bubble clknet_leaf_12_clk
+ sg13g2_dfrbpq_1
X_3373_ _1806_ net1003 _1805_ VPWR VGND sg13g2_nand2b_1
X_5112_ net1114 net1056 _0808_ VPWR VGND sg13g2_nor2b_1
X_6092_ net186 VGND VPWR _0142_ s0.data_out\[10\]\[7\] clknet_leaf_20_clk sg13g2_dfrbpq_2
X_5043_ s0.data_out\[15\]\[5\] s0.data_out\[14\]\[5\] net1133 _0748_ VPWR VGND sg13g2_mux2_1
XFILLER_26_727 VPWR VGND sg13g2_decap_8
XFILLER_26_749 VPWR VGND sg13g2_decap_8
X_5945_ VGND VPWR net1025 _1558_ _1559_ _1520_ sg13g2_a21oi_1
XFILLER_40_207 VPWR VGND sg13g2_decap_8
XFILLER_22_944 VPWR VGND sg13g2_fill_1
X_5876_ VGND VPWR _1496_ net487 net1328 sg13g2_or2_1
X_4827_ _0550_ net922 _0549_ VPWR VGND sg13g2_nand2_1
XFILLER_22_999 VPWR VGND sg13g2_decap_8
X_4758_ VPWR VGND _0422_ net1282 _0486_ net1275 _0487_ _0483_ sg13g2_a221oi_1
X_3709_ VGND VPWR _2108_ net576 net1309 sg13g2_or2_1
X_4689_ _0422_ _0425_ net1304 _0426_ VPWR VGND sg13g2_nand3_1
XFILLER_49_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_1017 VPWR VGND sg13g2_decap_8
XFILLER_0_336 VPWR VGND sg13g2_decap_8
XFILLER_1_837 VPWR VGND sg13g2_decap_8
XFILLER_0_369 VPWR VGND sg13g2_fill_1
XFILLER_29_510 VPWR VGND sg13g2_fill_2
XFILLER_29_521 VPWR VGND sg13g2_fill_2
XFILLER_1_1019 VPWR VGND sg13g2_decap_8
XFILLER_29_565 VPWR VGND sg13g2_fill_2
XFILLER_40_730 VPWR VGND sg13g2_decap_8
XFILLER_13_977 VPWR VGND sg13g2_decap_8
XFILLER_32_1010 VPWR VGND sg13g2_decap_8
XFILLER_4_631 VPWR VGND sg13g2_fill_1
XFILLER_4_620 VPWR VGND sg13g2_decap_4
XFILLER_4_686 VPWR VGND sg13g2_fill_1
XFILLER_4_697 VPWR VGND sg13g2_fill_2
Xhold3 s0.genblk1\[15\].modules.bubble VPWR VGND net299 sg13g2_dlygate4sd3_1
XFILLER_47_340 VPWR VGND sg13g2_decap_8
XFILLER_48_885 VPWR VGND sg13g2_decap_8
XFILLER_35_546 VPWR VGND sg13g2_fill_1
X_3991_ VGND VPWR _2364_ _2363_ _2314_ sg13g2_or2_1
X_5730_ _1363_ VPWR _1364_ VGND net1340 net428 sg13g2_o21ai_1
X_5661_ VPWR VGND _1240_ net1283 _1305_ net1278 _1306_ _1302_ sg13g2_a221oi_1
X_4612_ VGND VPWR _2825_ _0353_ _0354_ net1173 sg13g2_a21oi_1
X_5592_ _1244_ VPWR _1245_ VGND net1340 net404 sg13g2_o21ai_1
XFILLER_8_992 VPWR VGND sg13g2_decap_8
X_4543_ net1171 VPWR _0294_ VGND net1226 net1158 sg13g2_o21ai_1
X_4474_ net1170 net1049 _2792_ VPWR VGND sg13g2_nor2b_1
X_6213_ net175 VGND VPWR _0263_ s0.data_out\[0\]\[1\] clknet_leaf_7_clk sg13g2_dfrbpq_2
Xfanout916 _2469_ net916 VPWR VGND sg13g2_buf_8
X_3425_ net982 net1062 _1851_ VPWR VGND sg13g2_nor2b_1
X_3356_ _1788_ net995 _1763_ _1789_ VPWR VGND sg13g2_a21o_1
Xfanout927 _2460_ net927 VPWR VGND sg13g2_buf_1
Xfanout938 _2451_ net938 VPWR VGND sg13g2_buf_8
Xfanout949 net950 net949 VPWR VGND sg13g2_buf_2
X_6144_ net130 VGND VPWR _0194_ s0.data_out\[6\]\[4\] clknet_leaf_15_clk sg13g2_dfrbpq_2
X_6075_ net204 VGND VPWR _0125_ s0.data_out\[11\]\[2\] clknet_leaf_21_clk sg13g2_dfrbpq_2
X_3287_ _1726_ s0.data_out\[5\]\[2\] net1008 VPWR VGND sg13g2_nand2b_1
XFILLER_39_841 VPWR VGND sg13g2_fill_1
X_5026_ _0730_ net1123 _0702_ _0731_ VPWR VGND sg13g2_a21o_1
XFILLER_26_502 VPWR VGND sg13g2_fill_1
XFILLER_26_568 VPWR VGND sg13g2_fill_2
XFILLER_41_527 VPWR VGND sg13g2_fill_1
X_5928_ _1542_ net1023 _1541_ VPWR VGND sg13g2_nand2b_1
X_5859_ net1023 VPWR _1481_ VGND _1479_ _1480_ sg13g2_o21ai_1
XFILLER_10_947 VPWR VGND sg13g2_decap_8
X_6200__69 VPWR VGND net69 sg13g2_tiehi
XFILLER_1_634 VPWR VGND sg13g2_decap_8
XFILLER_0_144 VPWR VGND sg13g2_fill_2
XFILLER_0_122 VPWR VGND sg13g2_decap_8
XFILLER_0_199 VPWR VGND sg13g2_decap_8
XFILLER_29_340 VPWR VGND sg13g2_fill_2
XFILLER_45_844 VPWR VGND sg13g2_decap_8
XFILLER_29_395 VPWR VGND sg13g2_decap_8
XFILLER_40_571 VPWR VGND sg13g2_decap_8
XFILLER_9_723 VPWR VGND sg13g2_fill_2
XFILLER_8_244 VPWR VGND sg13g2_decap_8
XFILLER_8_288 VPWR VGND sg13g2_fill_2
XFILLER_5_951 VPWR VGND sg13g2_decap_8
XFILLER_4_483 VPWR VGND sg13g2_fill_2
X_4190_ net1190 s0.data_out\[20\]\[3\] _2535_ VPWR VGND sg13g2_and2_1
X_3210_ s0.data_out\[7\]\[1\] s0.data_out\[6\]\[1\] net1008 _1655_ VPWR VGND sg13g2_mux2_1
X_3141_ s0.data_out\[6\]\[0\] s0.data_out\[7\]\[0\] net1019 _1594_ VPWR VGND sg13g2_mux2_1
XFILLER_39_126 VPWR VGND sg13g2_fill_1
XFILLER_48_682 VPWR VGND sg13g2_decap_8
XFILLER_36_855 VPWR VGND sg13g2_decap_4
X_3974_ _2347_ net946 net345 VPWR VGND sg13g2_nand2_1
X_5713_ net1230 net1033 _1349_ VPWR VGND sg13g2_nor2b_1
XFILLER_31_560 VPWR VGND sg13g2_fill_2
X_5644_ net1039 net1047 _1290_ VPWR VGND sg13g2_nor2b_1
XFILLER_40_19 VPWR VGND sg13g2_decap_8
X_5575_ net1229 net1044 _1230_ VPWR VGND sg13g2_nor2b_1
Xhold211 s0.data_out\[13\]\[3\] VPWR VGND net507 sg13g2_dlygate4sd3_1
Xhold200 s0.data_out\[17\]\[1\] VPWR VGND net496 sg13g2_dlygate4sd3_1
Xhold222 _1649_ VPWR VGND net518 sg13g2_dlygate4sd3_1
Xhold233 _1019_ VPWR VGND net529 sg13g2_dlygate4sd3_1
X_4526_ s0.data_out\[19\]\[4\] s0.data_out\[18\]\[4\] net1176 _0279_ VPWR VGND sg13g2_mux2_1
Xhold244 s0.data_out\[11\]\[7\] VPWR VGND net540 sg13g2_dlygate4sd3_1
XFILLER_49_28 VPWR VGND sg13g2_decap_8
Xhold277 s0.data_out\[14\]\[2\] VPWR VGND net573 sg13g2_dlygate4sd3_1
Xhold255 s0.data_out\[19\]\[6\] VPWR VGND net551 sg13g2_dlygate4sd3_1
Xhold266 s0.data_out\[15\]\[6\] VPWR VGND net562 sg13g2_dlygate4sd3_1
X_4457_ _2777_ net927 _2776_ VPWR VGND sg13g2_nand2_1
Xhold299 s0.data_out\[8\]\[7\] VPWR VGND net595 sg13g2_dlygate4sd3_1
Xhold288 s0.data_out\[13\]\[7\] VPWR VGND net584 sg13g2_dlygate4sd3_1
X_3408_ net982 s0.data_out\[4\]\[1\] _1836_ VPWR VGND sg13g2_and2_1
X_6127_ net148 VGND VPWR _0177_ s0.valid_out\[7\][0] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_4388_ VGND VPWR net1197 _2715_ _2716_ _2676_ sg13g2_a21oi_1
X_3339_ VGND VPWR _1772_ _1771_ net1271 sg13g2_or2_1
X_6058_ net223 VGND VPWR _0108_ s0.genblk1\[12\].modules.bubble clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
XFILLER_22_1020 VPWR VGND sg13g2_decap_8
XFILLER_27_800 VPWR VGND sg13g2_fill_1
XFILLER_39_693 VPWR VGND sg13g2_fill_2
X_5009_ VGND VPWR net1122 _0713_ _0714_ _0661_ sg13g2_a21oi_1
XFILLER_42_825 VPWR VGND sg13g2_fill_2
XFILLER_6_704 VPWR VGND sg13g2_decap_8
XFILLER_10_755 VPWR VGND sg13g2_fill_1
XFILLER_5_269 VPWR VGND sg13g2_fill_2
XFILLER_5_247 VPWR VGND sg13g2_decap_4
XFILLER_30_63 VPWR VGND sg13g2_fill_1
XFILLER_30_74 VPWR VGND sg13g2_fill_1
XFILLER_2_910 VPWR VGND sg13g2_decap_8
XFILLER_2_987 VPWR VGND sg13g2_decap_8
XFILLER_1_475 VPWR VGND sg13g2_fill_1
XFILLER_49_457 VPWR VGND sg13g2_decap_8
XFILLER_39_61 VPWR VGND sg13g2_decap_4
XFILLER_29_181 VPWR VGND sg13g2_decap_8
XFILLER_17_354 VPWR VGND sg13g2_decap_4
XFILLER_18_888 VPWR VGND sg13g2_fill_2
XFILLER_44_173 VPWR VGND sg13g2_fill_2
XFILLER_18_899 VPWR VGND sg13g2_fill_2
XFILLER_41_891 VPWR VGND sg13g2_decap_8
XFILLER_9_586 VPWR VGND sg13g2_fill_1
X_3690_ net960 s0.data_out\[2\]\[4\] _2091_ VPWR VGND sg13g2_and2_1
X_5360_ VPWR _0114_ _1033_ VGND sg13g2_inv_1
X_4311_ _2645_ VPWR _2646_ VGND net1286 net455 sg13g2_o21ai_1
X_5291_ VGND VPWR net1118 _0971_ _0972_ _0931_ sg13g2_a21oi_1
X_4242_ VGND VPWR _2525_ _2576_ _2582_ net1273 sg13g2_a21oi_1
X_4173_ _0003_ _2516_ _2520_ _2482_ net1216 VPWR VGND sg13g2_a22oi_1
X_3124_ _1560_ _1562_ _1581_ VPWR VGND sg13g2_nor2b_1
XFILLER_28_619 VPWR VGND sg13g2_fill_1
XFILLER_23_335 VPWR VGND sg13g2_fill_2
X_3957_ VPWR _0255_ _2332_ VGND sg13g2_inv_1
XFILLER_13_1019 VPWR VGND sg13g2_decap_8
X_3888_ net1261 _2249_ _2273_ VPWR VGND sg13g2_nor2_1
X_5627_ _1275_ _2454_ _1274_ VPWR VGND sg13g2_nand2_1
X_5558_ s0.data_out\[11\]\[5\] s0.data_out\[10\]\[5\] net1085 _1215_ VPWR VGND sg13g2_mux2_1
X_4509_ _2825_ net1174 net579 VPWR VGND sg13g2_nand2_1
XFILLER_4_8 VPWR VGND sg13g2_fill_1
X_5489_ VGND VPWR _1151_ net486 net1335 sg13g2_or2_1
XFILLER_47_906 VPWR VGND sg13g2_decap_8
XFILLER_46_405 VPWR VGND sg13g2_decap_8
XFILLER_25_63 VPWR VGND sg13g2_fill_1
XFILLER_6_501 VPWR VGND sg13g2_fill_1
XFILLER_41_84 VPWR VGND sg13g2_decap_8
XFILLER_10_585 VPWR VGND sg13g2_decap_8
XFILLER_2_784 VPWR VGND sg13g2_decap_8
XFILLER_49_210 VPWR VGND sg13g2_decap_8
XFILLER_46_950 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_29_clk clknet_3_5__leaf_clk clknet_leaf_29_clk VPWR VGND sg13g2_buf_8
XFILLER_36_1008 VPWR VGND sg13g2_decap_8
X_4860_ net1136 net1051 _0579_ VPWR VGND sg13g2_nor2b_1
XFILLER_32_132 VPWR VGND sg13g2_fill_1
X_3811_ net961 VPWR _2201_ VGND _2199_ _2200_ sg13g2_o21ai_1
XFILLER_33_688 VPWR VGND sg13g2_fill_2
X_4791_ net1215 _0511_ _0516_ _0520_ VPWR VGND sg13g2_or3_1
X_3742_ VGND VPWR net973 _2138_ _2139_ _2111_ sg13g2_a21oi_1
X_3673_ _2076_ net932 _2075_ VPWR VGND sg13g2_nand2_1
X_5412_ _1028_ _1080_ _1081_ VPWR VGND sg13g2_and2_1
X_5343_ _1018_ VPWR _1019_ VGND _1014_ _1017_ sg13g2_o21ai_1
X_6135__140 VPWR VGND net140 sg13g2_tiehi
X_5274_ _0889_ VPWR _0955_ VGND net935 _0954_ sg13g2_o21ai_1
X_4225_ net364 net1207 _2566_ VPWR VGND sg13g2_nor2b_1
X_4156_ net1225 net1207 _2506_ VPWR VGND sg13g2_nor2b_1
X_3107_ _1564_ net1020 net411 VPWR VGND sg13g2_nand2_1
XFILLER_37_950 VPWR VGND sg13g2_decap_8
X_4087_ VPWR _2446_ net321 VGND sg13g2_inv_1
X_4989_ VGND VPWR net1125 s0.data_out\[14\]\[6\] _0696_ _0695_ sg13g2_a21oi_1
Xfanout1305 net1306 net1305 VPWR VGND sg13g2_buf_8
Xfanout1338 net1339 net1338 VPWR VGND sg13g2_buf_8
Xfanout1316 net1350 net1316 VPWR VGND sg13g2_buf_8
Xfanout1327 net1331 net1327 VPWR VGND sg13g2_buf_8
XFILLER_47_703 VPWR VGND sg13g2_decap_8
Xfanout1349 net1350 net1349 VPWR VGND sg13g2_buf_8
XFILLER_4_1028 VPWR VGND sg13g2_fill_1
XFILLER_28_961 VPWR VGND sg13g2_decap_4
XFILLER_36_95 VPWR VGND sg13g2_fill_1
XFILLER_15_622 VPWR VGND sg13g2_fill_2
XFILLER_27_493 VPWR VGND sg13g2_decap_4
XFILLER_43_975 VPWR VGND sg13g2_decap_8
XFILLER_15_655 VPWR VGND sg13g2_fill_1
XFILLER_42_474 VPWR VGND sg13g2_decap_8
XFILLER_30_658 VPWR VGND sg13g2_fill_1
XFILLER_10_371 VPWR VGND sg13g2_fill_1
X_6119__157 VPWR VGND net157 sg13g2_tiehi
XFILLER_2_581 VPWR VGND sg13g2_fill_2
XFILLER_2_570 VPWR VGND sg13g2_decap_8
X_4010_ VGND VPWR _2383_ _2382_ net1214 sg13g2_or2_1
XFILLER_28_4 VPWR VGND sg13g2_decap_4
XFILLER_38_725 VPWR VGND sg13g2_decap_4
XFILLER_37_202 VPWR VGND sg13g2_fill_1
XFILLER_37_235 VPWR VGND sg13g2_decap_8
X_5961_ net56 VGND VPWR _0011_ s0.shift_out\[21\][0] clknet_leaf_1_clk sg13g2_dfrbpq_2
XFILLER_19_994 VPWR VGND sg13g2_decap_8
XFILLER_45_290 VPWR VGND sg13g2_fill_1
X_4912_ _0629_ net1148 _0628_ VPWR VGND sg13g2_nand2b_1
XFILLER_34_942 VPWR VGND sg13g2_decap_8
X_5892_ _1506_ _1509_ net1330 _1510_ VPWR VGND sg13g2_nand3_1
X_4843_ _0564_ net923 _0563_ VPWR VGND sg13g2_nand2_1
XFILLER_21_614 VPWR VGND sg13g2_decap_8
XFILLER_21_625 VPWR VGND sg13g2_fill_2
XFILLER_21_647 VPWR VGND sg13g2_fill_1
X_4774_ VGND VPWR net1160 _0502_ _0503_ _0471_ sg13g2_a21oi_1
X_3725_ VGND VPWR net959 _2121_ _2122_ _2071_ sg13g2_a21oi_1
Xclkbuf_leaf_9_clk clknet_3_2__leaf_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
X_3656_ s0.data_out\[2\]\[0\] s0.data_out\[3\]\[0\] net976 _2061_ VPWR VGND sg13g2_mux2_1
X_3587_ net1309 VPWR _1997_ VGND net914 _1996_ sg13g2_o21ai_1
X_5326_ net1336 VPWR _1005_ VGND net408 _1000_ sg13g2_o21ai_1
X_5257_ net1107 net1048 _0939_ VPWR VGND sg13g2_nor2b_1
X_4208_ net1205 VPWR _2551_ VGND _2549_ _2550_ sg13g2_o21ai_1
X_5188_ net1229 net1110 _0879_ VPWR VGND sg13g2_nor2b_1
X_4139_ _2496_ VPWR net3 VGND _2481_ net913 sg13g2_o21ai_1
XFILLER_29_769 VPWR VGND sg13g2_decap_8
XFILLER_28_279 VPWR VGND sg13g2_fill_2
XFILLER_24_452 VPWR VGND sg13g2_fill_1
XFILLER_40_945 VPWR VGND sg13g2_decap_8
XFILLER_24_496 VPWR VGND sg13g2_fill_1
XFILLER_12_658 VPWR VGND sg13g2_fill_1
XFILLER_12_669 VPWR VGND sg13g2_decap_8
XFILLER_7_128 VPWR VGND sg13g2_decap_4
XFILLER_22_53 VPWR VGND sg13g2_fill_1
XFILLER_4_879 VPWR VGND sg13g2_decap_8
Xfanout1113 net1116 net1113 VPWR VGND sg13g2_buf_8
Xfanout1102 net1104 net1102 VPWR VGND sg13g2_buf_8
Xfanout1124 net1129 net1124 VPWR VGND sg13g2_buf_1
Xfanout1135 net1140 net1135 VPWR VGND sg13g2_buf_8
Xfanout1146 net1147 net1146 VPWR VGND sg13g2_buf_8
Xfanout1157 net1162 net1157 VPWR VGND sg13g2_buf_2
Xfanout1168 net1173 net1168 VPWR VGND sg13g2_buf_2
Xfanout1179 net1180 net1179 VPWR VGND sg13g2_buf_1
XFILLER_34_249 VPWR VGND sg13g2_decap_4
XFILLER_16_986 VPWR VGND sg13g2_decap_8
Xclkbuf_3_4__f_clk clknet_0_clk clknet_3_4__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_31_923 VPWR VGND sg13g2_fill_2
XFILLER_31_978 VPWR VGND sg13g2_decap_8
X_3510_ _1911_ _1912_ _1931_ VPWR VGND sg13g2_nor2b_1
X_4490_ VGND VPWR net1168 _2805_ _2806_ _2765_ sg13g2_a21oi_1
X_3441_ net984 net1054 _1865_ VPWR VGND sg13g2_nor2b_1
X_6160_ net113 VGND VPWR _0210_ s0.shift_out\[5\][0] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_3372_ VGND VPWR net992 _1804_ _1805_ _1743_ sg13g2_a21oi_1
X_5111_ VGND VPWR _0747_ _0806_ _0807_ net1128 sg13g2_a21oi_1
X_6091_ net187 VGND VPWR _0141_ s0.data_out\[10\]\[6\] clknet_leaf_20_clk sg13g2_dfrbpq_2
X_6132__143 VPWR VGND net143 sg13g2_tiehi
X_5042_ _0747_ net1132 net548 VPWR VGND sg13g2_nand2_1
XFILLER_19_0 VPWR VGND sg13g2_fill_1
XFILLER_38_566 VPWR VGND sg13g2_fill_2
X_5944_ _1557_ net1017 _1521_ _1558_ VPWR VGND sg13g2_a21o_1
X_5875_ net1328 VPWR _1495_ VGND net918 _1494_ sg13g2_o21ai_1
X_4826_ s0.data_out\[15\]\[2\] s0.data_out\[16\]\[2\] net1152 _0549_ VPWR VGND sg13g2_mux2_1
XFILLER_21_444 VPWR VGND sg13g2_decap_8
XFILLER_22_978 VPWR VGND sg13g2_decap_8
X_4757_ _0486_ net1160 _0485_ VPWR VGND sg13g2_nand2b_1
X_3708_ net1309 VPWR _2107_ VGND net933 _2106_ sg13g2_o21ai_1
X_4688_ net1160 VPWR _0425_ VGND _0423_ _0424_ sg13g2_o21ai_1
X_3639_ VGND VPWR _2031_ _2046_ _2048_ _1937_ sg13g2_a21oi_1
XFILLER_1_816 VPWR VGND sg13g2_decap_8
XFILLER_0_315 VPWR VGND sg13g2_decap_8
X_5309_ _0990_ net1215 _0981_ VPWR VGND sg13g2_xnor2_1
XFILLER_29_533 VPWR VGND sg13g2_decap_8
XFILLER_29_577 VPWR VGND sg13g2_fill_2
XFILLER_44_547 VPWR VGND sg13g2_fill_1
XFILLER_44_536 VPWR VGND sg13g2_decap_4
XFILLER_17_75 VPWR VGND sg13g2_decap_8
XFILLER_13_912 VPWR VGND sg13g2_fill_1
XFILLER_13_956 VPWR VGND sg13g2_decap_8
XFILLER_40_786 VPWR VGND sg13g2_decap_8
XFILLER_8_437 VPWR VGND sg13g2_fill_2
X_5962__55 VPWR VGND net55 sg13g2_tiehi
X_6079__200 VPWR VGND net200 sg13g2_tiehi
XFILLER_3_175 VPWR VGND sg13g2_fill_1
Xhold4 s0.genblk1\[2\].modules.bubble VPWR VGND net300 sg13g2_dlygate4sd3_1
XFILLER_48_864 VPWR VGND sg13g2_decap_8
XFILLER_47_330 VPWR VGND sg13g2_decap_4
XFILLER_35_514 VPWR VGND sg13g2_fill_2
X_3990_ VGND VPWR _2361_ _2362_ _2363_ _2465_ sg13g2_a21oi_1
XFILLER_15_260 VPWR VGND sg13g2_decap_8
XFILLER_43_591 VPWR VGND sg13g2_fill_1
X_5660_ _1305_ net1078 _1304_ VPWR VGND sg13g2_nand2b_1
XFILLER_30_230 VPWR VGND sg13g2_fill_1
X_4611_ _0353_ net341 net1175 VPWR VGND sg13g2_nand2b_1
XFILLER_30_241 VPWR VGND sg13g2_fill_1
XFILLER_30_252 VPWR VGND sg13g2_fill_2
X_5591_ _1240_ _1243_ net1340 _1244_ VPWR VGND sg13g2_nand3_1
XFILLER_30_296 VPWR VGND sg13g2_fill_2
XFILLER_8_971 VPWR VGND sg13g2_decap_8
X_4542_ net1303 net304 _0036_ VPWR VGND sg13g2_and2_1
XFILLER_7_492 VPWR VGND sg13g2_fill_1
X_4473_ VGND VPWR _2713_ _2790_ _2791_ net1184 sg13g2_a21oi_1
X_6212_ net195 VGND VPWR _0262_ s0.data_out\[0\]\[0\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_3424_ net982 s0.data_out\[4\]\[3\] _1850_ VPWR VGND sg13g2_and2_1
X_3355_ s0.data_out\[6\]\[7\] s0.data_out\[5\]\[7\] net998 _1788_ VPWR VGND sg13g2_mux2_1
Xfanout928 _2459_ net928 VPWR VGND sg13g2_buf_8
Xfanout939 _2448_ net939 VPWR VGND sg13g2_buf_8
X_6143_ net131 VGND VPWR _0193_ s0.data_out\[6\]\[3\] clknet_leaf_15_clk sg13g2_dfrbpq_2
Xfanout917 _2468_ net917 VPWR VGND sg13g2_buf_8
X_6074_ net205 VGND VPWR _0124_ s0.data_out\[11\]\[1\] clknet_leaf_25_clk sg13g2_dfrbpq_2
X_3286_ VPWR _0191_ _1725_ VGND sg13g2_inv_1
XFILLER_38_330 VPWR VGND sg13g2_decap_4
X_5025_ s0.data_out\[15\]\[7\] s0.data_out\[14\]\[7\] net1130 _0730_ VPWR VGND sg13g2_mux2_1
XFILLER_0_1020 VPWR VGND sg13g2_decap_8
X_5927_ VGND VPWR net1013 _1540_ _1541_ _1480_ sg13g2_a21oi_1
XFILLER_34_591 VPWR VGND sg13g2_decap_8
XFILLER_10_926 VPWR VGND sg13g2_decap_8
XFILLER_16_1028 VPWR VGND sg13g2_fill_1
XFILLER_22_764 VPWR VGND sg13g2_decap_4
X_5858_ net1013 net1075 _1480_ VPWR VGND sg13g2_nor2b_1
XFILLER_6_919 VPWR VGND sg13g2_decap_8
X_4809_ net1220 _0527_ _0528_ _0062_ VPWR VGND sg13g2_nor3_1
X_5789_ _1414_ VPWR _1415_ VGND net1031 _2489_ sg13g2_o21ai_1
XFILLER_1_613 VPWR VGND sg13g2_decap_8
XFILLER_49_639 VPWR VGND sg13g2_decap_8
XFILLER_0_178 VPWR VGND sg13g2_decap_8
XFILLER_45_823 VPWR VGND sg13g2_decap_8
XFILLER_44_311 VPWR VGND sg13g2_fill_2
XFILLER_28_85 VPWR VGND sg13g2_fill_1
XFILLER_44_355 VPWR VGND sg13g2_fill_1
XFILLER_9_757 VPWR VGND sg13g2_decap_4
XFILLER_12_296 VPWR VGND sg13g2_decap_8
XFILLER_5_930 VPWR VGND sg13g2_decap_8
X_3140_ net1220 _1586_ _1591_ _0177_ VPWR VGND sg13g2_nor3_1
XFILLER_48_661 VPWR VGND sg13g2_decap_8
XFILLER_36_801 VPWR VGND sg13g2_decap_8
XFILLER_10_4 VPWR VGND sg13g2_fill_1
XFILLER_36_834 VPWR VGND sg13g2_fill_1
XFILLER_39_1028 VPWR VGND sg13g2_fill_1
XFILLER_23_539 VPWR VGND sg13g2_fill_1
X_3973_ VPWR _0257_ _2346_ VGND sg13g2_inv_1
X_5712_ net1037 VPWR _1348_ VGND net1230 net1028 sg13g2_o21ai_1
X_5643_ VGND VPWR _1199_ _1288_ _1289_ net1083 sg13g2_a21oi_1
X_5574_ net1082 VPWR _1229_ VGND net1229 net1039 sg13g2_o21ai_1
Xhold201 _0434_ VPWR VGND net497 sg13g2_dlygate4sd3_1
X_4525_ _0278_ net1248 _0277_ VPWR VGND sg13g2_nand2_1
Xhold223 s0.data_out\[6\]\[7\] VPWR VGND net519 sg13g2_dlygate4sd3_1
Xhold212 _0915_ VPWR VGND net508 sg13g2_dlygate4sd3_1
Xhold234 s0.data_out\[17\]\[2\] VPWR VGND net530 sg13g2_dlygate4sd3_1
Xhold278 s0.data_out\[19\]\[7\] VPWR VGND net574 sg13g2_dlygate4sd3_1
Xhold256 _2796_ VPWR VGND net552 sg13g2_dlygate4sd3_1
Xhold267 _0699_ VPWR VGND net563 sg13g2_dlygate4sd3_1
X_4456_ s0.data_out\[18\]\[4\] s0.data_out\[19\]\[4\] net1188 _2776_ VPWR VGND sg13g2_mux2_1
Xhold245 s0.data_out\[11\]\[5\] VPWR VGND net541 sg13g2_dlygate4sd3_1
Xhold289 _0943_ VPWR VGND net585 sg13g2_dlygate4sd3_1
X_4387_ _2714_ net1182 _2677_ _2715_ VPWR VGND sg13g2_a21o_1
X_3407_ _1835_ net915 _1834_ VPWR VGND sg13g2_nand2_1
X_6126_ net150 VGND VPWR net327 s0.was_valid_out\[7\][0] clknet_leaf_16_clk sg13g2_dfrbpq_2
X_3338_ VGND VPWR net1000 _1770_ _1771_ _1727_ sg13g2_a21oi_1
X_3269_ _1710_ _1711_ _0188_ VPWR VGND sg13g2_nor2_1
X_6057_ net224 VGND VPWR _0107_ s0.shift_out\[13\][0] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_5008_ s0.data_out\[15\]\[1\] s0.data_out\[14\]\[1\] net1130 _0713_ VPWR VGND sg13g2_mux2_1
XFILLER_26_311 VPWR VGND sg13g2_fill_2
XFILLER_42_859 VPWR VGND sg13g2_decap_8
XFILLER_10_778 VPWR VGND sg13g2_fill_2
XFILLER_5_215 VPWR VGND sg13g2_fill_1
X_6076__203 VPWR VGND net203 sg13g2_tiehi
XFILLER_30_53 VPWR VGND sg13g2_fill_1
XFILLER_2_966 VPWR VGND sg13g2_decap_8
XFILLER_1_443 VPWR VGND sg13g2_decap_4
XFILLER_49_436 VPWR VGND sg13g2_decap_8
XFILLER_44_141 VPWR VGND sg13g2_fill_2
XFILLER_18_867 VPWR VGND sg13g2_decap_8
XFILLER_45_697 VPWR VGND sg13g2_decap_8
XFILLER_45_675 VPWR VGND sg13g2_decap_8
XFILLER_17_399 VPWR VGND sg13g2_decap_4
XFILLER_9_598 VPWR VGND sg13g2_fill_1
XFILLER_5_782 VPWR VGND sg13g2_fill_1
X_4310_ _2641_ _2644_ net1286 _2645_ VPWR VGND sg13g2_nand3_1
X_5290_ _0970_ net1107 _0932_ _0971_ VPWR VGND sg13g2_a21o_1
XFILLER_4_292 VPWR VGND sg13g2_fill_2
X_4241_ net1281 _2580_ _2581_ VPWR VGND sg13g2_nor2_1
X_4172_ net1216 _2519_ _2520_ VPWR VGND sg13g2_nor2_1
X_3123_ _1563_ _1579_ _1580_ VPWR VGND sg13g2_nor2b_1
XFILLER_27_119 VPWR VGND sg13g2_fill_2
X_3956_ _2331_ VPWR _2332_ VGND net1295 net479 sg13g2_o21ai_1
XFILLER_11_509 VPWR VGND sg13g2_decap_8
X_3887_ _2212_ _2271_ net1247 _2272_ VPWR VGND sg13g2_nand3_1
X_5626_ _1214_ VPWR _1274_ VGND net1087 _2490_ sg13g2_o21ai_1
XFILLER_31_391 VPWR VGND sg13g2_fill_1
X_5557_ _1214_ net1086 s0.data_out\[10\]\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_3_719 VPWR VGND sg13g2_decap_8
X_4508_ _2818_ _2823_ _2824_ VPWR VGND sg13g2_nor2_1
XFILLER_2_207 VPWR VGND sg13g2_fill_2
X_5488_ net1335 VPWR _1150_ VGND net939 _1149_ sg13g2_o21ai_1
X_4439_ VPWR _0028_ _2761_ VGND sg13g2_inv_1
X_6109_ net168 VGND VPWR _0159_ s0.data_out\[9\]\[5\] clknet_leaf_18_clk sg13g2_dfrbpq_2
XFILLER_26_185 VPWR VGND sg13g2_decap_4
XFILLER_10_542 VPWR VGND sg13g2_fill_1
XFILLER_29_1016 VPWR VGND sg13g2_decap_8
XFILLER_29_1027 VPWR VGND sg13g2_fill_2
XFILLER_2_763 VPWR VGND sg13g2_decap_8
XFILLER_1_284 VPWR VGND sg13g2_fill_2
XFILLER_49_266 VPWR VGND sg13g2_decap_4
XFILLER_37_406 VPWR VGND sg13g2_fill_2
X_5987__28 VPWR VGND net28 sg13g2_tiehi
XFILLER_45_483 VPWR VGND sg13g2_fill_1
XFILLER_33_645 VPWR VGND sg13g2_fill_2
X_4790_ _0508_ _0516_ _0517_ _0518_ _0519_ VPWR VGND sg13g2_nor4_1
X_3810_ net950 net1061 _2200_ VPWR VGND sg13g2_nor2b_1
X_3741_ _2137_ net963 _2112_ _2138_ VPWR VGND sg13g2_a21o_1
XFILLER_32_188 VPWR VGND sg13g2_decap_4
XFILLER_12_1020 VPWR VGND sg13g2_decap_8
X_3672_ s0.data_out\[2\]\[2\] s0.data_out\[3\]\[2\] net976 _2075_ VPWR VGND sg13g2_mux2_1
X_5411_ _1080_ net1103 _1079_ VPWR VGND sg13g2_nand2b_1
X_5342_ VGND VPWR _1018_ net528 net1334 sg13g2_or2_1
XFILLER_49_0 VPWR VGND sg13g2_decap_8
X_5273_ VGND VPWR net1100 _0953_ _0954_ _0891_ sg13g2_a21oi_1
X_4224_ net1203 VPWR _2565_ VGND _2563_ _2564_ sg13g2_o21ai_1
X_4155_ VGND VPWR _2505_ _2504_ _2503_ sg13g2_or2_1
XFILLER_28_439 VPWR VGND sg13g2_fill_2
X_4086_ VPWR _2445_ net346 VGND sg13g2_inv_1
X_4988_ net1125 net1051 _0695_ VPWR VGND sg13g2_nor2b_1
X_3939_ VGND VPWR _2317_ net513 net1293 sg13g2_or2_1
XFILLER_20_884 VPWR VGND sg13g2_fill_1
X_5609_ VPWR _0137_ _1259_ VGND sg13g2_inv_1
XFILLER_3_516 VPWR VGND sg13g2_fill_1
X_6073__206 VPWR VGND net206 sg13g2_tiehi
Xfanout1317 net1318 net1317 VPWR VGND sg13g2_buf_8
Xfanout1306 net1316 net1306 VPWR VGND sg13g2_buf_8
Xfanout1339 net1349 net1339 VPWR VGND sg13g2_buf_8
Xfanout1328 net1331 net1328 VPWR VGND sg13g2_buf_2
XFILLER_46_214 VPWR VGND sg13g2_decap_4
XFILLER_46_203 VPWR VGND sg13g2_fill_2
XFILLER_47_759 VPWR VGND sg13g2_decap_8
XFILLER_27_461 VPWR VGND sg13g2_decap_4
XFILLER_43_954 VPWR VGND sg13g2_decap_8
XFILLER_42_431 VPWR VGND sg13g2_fill_1
XFILLER_15_678 VPWR VGND sg13g2_fill_2
XFILLER_35_1020 VPWR VGND sg13g2_decap_8
XFILLER_15_689 VPWR VGND sg13g2_fill_2
XFILLER_14_199 VPWR VGND sg13g2_fill_1
XFILLER_42_7 VPWR VGND sg13g2_fill_2
XFILLER_42_1013 VPWR VGND sg13g2_decap_8
XFILLER_38_748 VPWR VGND sg13g2_fill_1
XFILLER_38_715 VPWR VGND sg13g2_fill_1
XFILLER_37_214 VPWR VGND sg13g2_decap_8
X_5960_ net57 VGND VPWR net365 s0.data_out\[21\]\[7\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_19_973 VPWR VGND sg13g2_decap_8
X_5891_ net1025 VPWR _1509_ VGND _1507_ _1508_ sg13g2_o21ai_1
X_4911_ VGND VPWR net1136 _0627_ _0628_ _0566_ sg13g2_a21oi_1
XFILLER_33_442 VPWR VGND sg13g2_fill_1
X_4842_ s0.data_out\[15\]\[4\] s0.data_out\[16\]\[4\] net1153 _0563_ VPWR VGND sg13g2_mux2_1
XFILLER_34_998 VPWR VGND sg13g2_decap_8
X_4773_ _0501_ net1145 _0472_ _0502_ VPWR VGND sg13g2_a21o_1
X_3724_ s0.data_out\[3\]\[1\] s0.data_out\[2\]\[1\] net965 _2121_ VPWR VGND sg13g2_mux2_1
X_3655_ net1219 _2055_ _0225_ VPWR VGND sg13g2_nor2_1
X_3586_ VGND VPWR net972 net515 _1996_ _1995_ sg13g2_a21oi_1
X_5325_ VGND VPWR _0998_ _1001_ _1004_ _1003_ sg13g2_a21oi_1
X_5256_ VGND VPWR _0846_ _0937_ _0938_ net1118 sg13g2_a21oi_1
X_4207_ net1195 net1053 _2550_ VPWR VGND sg13g2_nor2b_1
X_5187_ net1117 VPWR _0878_ VGND net1229 net1106 sg13g2_o21ai_1
X_4138_ _2496_ net1273 net913 VPWR VGND sg13g2_nand2_1
X_4069_ net1274 _2402_ _2403_ _2430_ VPWR VGND sg13g2_nor3_1
XFILLER_19_1015 VPWR VGND sg13g2_decap_8
X_5974__42 VPWR VGND net42 sg13g2_tiehi
XFILLER_24_475 VPWR VGND sg13g2_decap_4
XFILLER_8_619 VPWR VGND sg13g2_decap_8
XFILLER_11_147 VPWR VGND sg13g2_fill_1
XFILLER_22_43 VPWR VGND sg13g2_fill_1
XFILLER_22_65 VPWR VGND sg13g2_fill_2
XFILLER_4_858 VPWR VGND sg13g2_decap_8
XFILLER_3_335 VPWR VGND sg13g2_decap_8
XFILLER_3_313 VPWR VGND sg13g2_fill_2
Xfanout1103 net1104 net1103 VPWR VGND sg13g2_buf_1
XFILLER_26_1008 VPWR VGND sg13g2_decap_8
Xfanout1114 net1116 net1114 VPWR VGND sg13g2_buf_8
Xfanout1125 net1129 net1125 VPWR VGND sg13g2_buf_8
Xfanout1147 net1150 net1147 VPWR VGND sg13g2_buf_8
Xfanout1136 net1137 net1136 VPWR VGND sg13g2_buf_8
Xfanout1169 net1173 net1169 VPWR VGND sg13g2_buf_8
Xfanout1158 net1159 net1158 VPWR VGND sg13g2_buf_8
XFILLER_47_534 VPWR VGND sg13g2_decap_4
XFILLER_47_62 VPWR VGND sg13g2_fill_1
XFILLER_47_589 VPWR VGND sg13g2_fill_2
XFILLER_47_578 VPWR VGND sg13g2_decap_8
XFILLER_27_291 VPWR VGND sg13g2_fill_1
XFILLER_43_784 VPWR VGND sg13g2_fill_1
XFILLER_42_250 VPWR VGND sg13g2_decap_4
XFILLER_31_935 VPWR VGND sg13g2_decap_8
XFILLER_31_946 VPWR VGND sg13g2_fill_1
X_6125__151 VPWR VGND net151 sg13g2_tiehi
XFILLER_30_456 VPWR VGND sg13g2_fill_2
XFILLER_31_957 VPWR VGND sg13g2_decap_8
X_3440_ net984 s0.data_out\[4\]\[5\] _1864_ VPWR VGND sg13g2_and2_1
X_3371_ s0.data_out\[6\]\[4\] s0.data_out\[5\]\[4\] net999 _1804_ VPWR VGND sg13g2_mux2_1
X_6090_ net188 VGND VPWR _0140_ s0.data_out\[10\]\[5\] clknet_leaf_19_clk sg13g2_dfrbpq_2
XFILLER_3_880 VPWR VGND sg13g2_decap_8
X_5110_ _0806_ s0.data_out\[13\]\[5\] net1132 VPWR VGND sg13g2_nand2b_1
X_5041_ VGND VPWR _0746_ _0745_ net1215 sg13g2_or2_1
XFILLER_26_707 VPWR VGND sg13g2_fill_1
X_5943_ s0.data_out\[8\]\[6\] s0.data_out\[7\]\[6\] net1021 _1557_ VPWR VGND sg13g2_mux2_1
XFILLER_21_412 VPWR VGND sg13g2_decap_8
XFILLER_22_935 VPWR VGND sg13g2_decap_8
X_5874_ VGND VPWR net1013 net467 _1494_ _1493_ sg13g2_a21oi_1
XFILLER_33_261 VPWR VGND sg13g2_fill_2
X_4825_ VPWR _0064_ _0548_ VGND sg13g2_inv_1
XFILLER_22_957 VPWR VGND sg13g2_fill_2
X_5971__45 VPWR VGND net45 sg13g2_tiehi
X_4756_ VGND VPWR net1144 _0484_ _0485_ _0424_ sg13g2_a21oi_1
X_3707_ VGND VPWR net964 net491 _2106_ _2105_ sg13g2_a21oi_1
X_4687_ net1144 net1073 _0424_ VPWR VGND sg13g2_nor2b_1
X_3638_ _2047_ _2030_ _2028_ VPWR VGND sg13g2_nand2b_1
X_3569_ net972 s0.data_out\[3\]\[5\] _1981_ VPWR VGND sg13g2_and2_1
X_5308_ net1265 _0961_ _0989_ VPWR VGND sg13g2_nor2_1
X_5239_ _0923_ net501 net1121 VPWR VGND sg13g2_nand2b_1
XFILLER_29_523 VPWR VGND sg13g2_fill_1
XFILLER_17_707 VPWR VGND sg13g2_decap_8
XFILLER_25_740 VPWR VGND sg13g2_decap_8
XFILLER_13_935 VPWR VGND sg13g2_decap_8
X_6109__168 VPWR VGND net168 sg13g2_tiehi
XFILLER_21_990 VPWR VGND sg13g2_decap_8
XFILLER_4_655 VPWR VGND sg13g2_fill_2
XFILLER_4_699 VPWR VGND sg13g2_fill_1
XFILLER_48_843 VPWR VGND sg13g2_decap_8
XFILLER_0_894 VPWR VGND sg13g2_decap_8
XFILLER_12_8 VPWR VGND sg13g2_fill_2
Xhold5 s0.genblk1\[20\].modules.bubble VPWR VGND net301 sg13g2_dlygate4sd3_1
XFILLER_16_773 VPWR VGND sg13g2_decap_8
XFILLER_31_732 VPWR VGND sg13g2_decap_8
X_4610_ VPWR _0045_ net559 VGND sg13g2_inv_1
XFILLER_31_776 VPWR VGND sg13g2_fill_1
XFILLER_8_950 VPWR VGND sg13g2_decap_8
X_5590_ net1077 VPWR _1243_ VGND _1241_ _1242_ sg13g2_o21ai_1
X_4541_ VGND VPWR _0288_ _0292_ _0035_ _0293_ sg13g2_a21oi_1
X_4472_ _2790_ s0.data_out\[18\]\[6\] net1189 VPWR VGND sg13g2_nand2b_1
X_6211_ net208 VGND VPWR _0261_ s0.valid_out\[0\][0] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_3423_ _1849_ net915 _1848_ VPWR VGND sg13g2_nand2_1
X_6142_ net132 VGND VPWR _0192_ s0.data_out\[6\]\[2\] clknet_leaf_15_clk sg13g2_dfrbpq_2
X_3354_ _1787_ net998 net569 VPWR VGND sg13g2_nand2_1
Xfanout918 _2467_ net918 VPWR VGND sg13g2_buf_8
Xfanout929 _2459_ net929 VPWR VGND sg13g2_buf_1
XFILLER_31_0 VPWR VGND sg13g2_decap_4
X_6073_ net206 VGND VPWR _0123_ s0.data_out\[11\]\[0\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_3285_ _1724_ VPWR _1725_ VGND _1720_ _1723_ sg13g2_o21ai_1
XFILLER_39_832 VPWR VGND sg13g2_fill_2
X_5024_ _0729_ net1131 net577 VPWR VGND sg13g2_nand2_1
XFILLER_38_397 VPWR VGND sg13g2_fill_1
XFILLER_26_515 VPWR VGND sg13g2_decap_4
XFILLER_0_90 VPWR VGND sg13g2_fill_2
X_5926_ s0.data_out\[8\]\[0\] s0.data_out\[7\]\[0\] net1019 _1540_ VPWR VGND sg13g2_mux2_1
XFILLER_16_1007 VPWR VGND sg13g2_decap_8
X_5857_ net1012 s0.data_out\[7\]\[0\] _1479_ VPWR VGND sg13g2_and2_1
X_4808_ VGND VPWR _2446_ _0529_ _0061_ _0534_ sg13g2_a21oi_1
X_5788_ _1414_ net1031 net487 VPWR VGND sg13g2_nand2_1
XFILLER_5_408 VPWR VGND sg13g2_decap_4
X_4739_ VPWR _0057_ _0469_ VGND sg13g2_inv_1
XFILLER_1_669 VPWR VGND sg13g2_decap_8
XFILLER_49_618 VPWR VGND sg13g2_decap_8
X_6115__161 VPWR VGND net161 sg13g2_tiehi
XFILLER_45_802 VPWR VGND sg13g2_decap_8
XFILLER_44_323 VPWR VGND sg13g2_fill_2
XFILLER_29_375 VPWR VGND sg13g2_fill_2
XFILLER_45_879 VPWR VGND sg13g2_decap_8
XFILLER_8_213 VPWR VGND sg13g2_decap_8
X_6122__154 VPWR VGND net154 sg13g2_tiehi
XFILLER_5_986 VPWR VGND sg13g2_decap_8
XFILLER_4_485 VPWR VGND sg13g2_fill_1
XFILLER_0_691 VPWR VGND sg13g2_decap_8
XFILLER_48_640 VPWR VGND sg13g2_decap_8
XFILLER_39_1007 VPWR VGND sg13g2_decap_8
X_3972_ _2345_ VPWR _2346_ VGND _2341_ _2344_ sg13g2_o21ai_1
XFILLER_16_592 VPWR VGND sg13g2_fill_2
X_5711_ net1045 net1231 net1223 _0151_ VPWR VGND sg13g2_mux2_1
X_5642_ _1288_ s0.data_out\[9\]\[7\] net1086 VPWR VGND sg13g2_nand2b_1
X_5573_ net1346 net315 _0132_ VPWR VGND sg13g2_and2_1
XFILLER_8_791 VPWR VGND sg13g2_fill_2
Xhold202 s0.data_out\[18\]\[2\] VPWR VGND net498 sg13g2_dlygate4sd3_1
X_4524_ VGND VPWR net1184 _0276_ _0277_ _2784_ sg13g2_a21oi_1
Xhold224 _1767_ VPWR VGND net520 sg13g2_dlygate4sd3_1
Xhold213 s0.data_out\[3\]\[3\] VPWR VGND net509 sg13g2_dlygate4sd3_1
Xhold235 s0.data_out\[10\]\[7\] VPWR VGND net531 sg13g2_dlygate4sd3_1
Xhold257 s0.data_out\[2\]\[7\] VPWR VGND net553 sg13g2_dlygate4sd3_1
Xhold246 s0.data_out\[9\]\[6\] VPWR VGND net542 sg13g2_dlygate4sd3_1
X_4455_ VPWR _0030_ _2775_ VGND sg13g2_inv_1
Xhold268 s0.data_out\[14\]\[1\] VPWR VGND net564 sg13g2_dlygate4sd3_1
Xhold279 _2803_ VPWR VGND net575 sg13g2_dlygate4sd3_1
X_4386_ s0.data_out\[20\]\[6\] s0.data_out\[19\]\[6\] net1188 _2714_ VPWR VGND sg13g2_mux2_1
X_3406_ s0.data_out\[4\]\[1\] s0.data_out\[5\]\[1\] net997 _1834_ VPWR VGND sg13g2_mux2_1
X_6125_ net151 VGND VPWR _0175_ s0.genblk1\[7\].modules.bubble clknet_leaf_17_clk
+ sg13g2_dfrbpq_1
X_3337_ _1769_ net991 _1728_ _1770_ VPWR VGND sg13g2_a21o_1
X_3268_ net1325 VPWR _1711_ VGND net465 _1706_ sg13g2_o21ai_1
X_6056_ net225 VGND VPWR _0106_ s0.data_out\[13\]\[7\] clknet_leaf_27_clk sg13g2_dfrbpq_2
X_3199_ net1006 net1047 _1645_ VPWR VGND sg13g2_nor2b_1
XFILLER_38_150 VPWR VGND sg13g2_decap_4
X_5007_ _0712_ net1131 net564 VPWR VGND sg13g2_nand2_1
X_6069__211 VPWR VGND net211 sg13g2_tiehi
XFILLER_27_813 VPWR VGND sg13g2_decap_4
XFILLER_27_835 VPWR VGND sg13g2_decap_4
X_5909_ _1524_ VPWR _1525_ VGND _1520_ _1523_ sg13g2_o21ai_1
XFILLER_30_21 VPWR VGND sg13g2_decap_8
XFILLER_30_32 VPWR VGND sg13g2_fill_1
XFILLER_2_945 VPWR VGND sg13g2_decap_8
XFILLER_49_415 VPWR VGND sg13g2_decap_8
XFILLER_7_1027 VPWR VGND sg13g2_fill_2
XFILLER_18_813 VPWR VGND sg13g2_fill_2
XFILLER_44_186 VPWR VGND sg13g2_fill_2
XFILLER_44_175 VPWR VGND sg13g2_fill_1
XFILLER_9_566 VPWR VGND sg13g2_fill_2
XFILLER_9_577 VPWR VGND sg13g2_decap_8
XFILLER_5_750 VPWR VGND sg13g2_fill_2
X_4240_ VGND VPWR net1202 _2579_ _2580_ _2519_ sg13g2_a21oi_1
X_4171_ net1202 _2517_ _2518_ _2519_ VPWR VGND sg13g2_nor3_1
X_3122_ _1573_ VPWR _1579_ VGND _1568_ _1575_ sg13g2_o21ai_1
XFILLER_49_982 VPWR VGND sg13g2_decap_8
XFILLER_48_492 VPWR VGND sg13g2_decap_8
X_3955_ _2327_ _2330_ net1295 _2331_ VPWR VGND sg13g2_nand3_1
X_3886_ _2271_ net962 _2270_ VPWR VGND sg13g2_nand2b_1
X_5625_ VPWR _0139_ _1273_ VGND sg13g2_inv_1
X_5556_ VGND VPWR net1093 _1212_ _1213_ _1154_ sg13g2_a21oi_1
X_4507_ _2822_ VPWR _2823_ VGND net1212 _2807_ sg13g2_o21ai_1
X_5487_ VGND VPWR net1078 net436 _1149_ _1148_ sg13g2_a21oi_1
X_4438_ _2760_ VPWR _2761_ VGND net1287 net464 sg13g2_o21ai_1
X_4369_ _2641_ _2696_ _2697_ VPWR VGND sg13g2_and2_1
X_6108_ net169 VGND VPWR _0158_ s0.data_out\[9\]\[4\] clknet_leaf_19_clk sg13g2_dfrbpq_2
XFILLER_46_418 VPWR VGND sg13g2_decap_4
X_6039_ net243 VGND VPWR _0089_ s0.data_out\[14\]\[2\] clknet_leaf_29_clk sg13g2_dfrbpq_2
XFILLER_27_643 VPWR VGND sg13g2_decap_8
XFILLER_27_676 VPWR VGND sg13g2_fill_2
XFILLER_25_32 VPWR VGND sg13g2_fill_2
XFILLER_42_657 VPWR VGND sg13g2_fill_1
XFILLER_41_156 VPWR VGND sg13g2_fill_2
XFILLER_41_145 VPWR VGND sg13g2_fill_1
XFILLER_30_808 VPWR VGND sg13g2_decap_8
XFILLER_30_819 VPWR VGND sg13g2_fill_1
XFILLER_23_871 VPWR VGND sg13g2_decap_8
XFILLER_10_521 VPWR VGND sg13g2_decap_8
XFILLER_6_514 VPWR VGND sg13g2_decap_8
XFILLER_6_558 VPWR VGND sg13g2_fill_2
XFILLER_2_742 VPWR VGND sg13g2_decap_8
XFILLER_49_234 VPWR VGND sg13g2_decap_8
XFILLER_38_919 VPWR VGND sg13g2_decap_8
XFILLER_37_418 VPWR VGND sg13g2_fill_1
XFILLER_46_985 VPWR VGND sg13g2_decap_8
XFILLER_17_197 VPWR VGND sg13g2_decap_8
XFILLER_33_668 VPWR VGND sg13g2_decap_8
X_3740_ s0.data_out\[3\]\[7\] s0.data_out\[2\]\[7\] net967 _2137_ VPWR VGND sg13g2_mux2_1
X_3671_ VPWR _0227_ _2074_ VGND sg13g2_inv_1
XFILLER_9_396 VPWR VGND sg13g2_fill_2
X_5410_ VGND VPWR net1089 _1078_ _1079_ _1030_ sg13g2_a21oi_1
X_5341_ net1334 VPWR _1017_ VGND net938 _1016_ sg13g2_o21ai_1
X_5272_ s0.data_out\[13\]\[0\] s0.data_out\[12\]\[0\] net1108 _0953_ VPWR VGND sg13g2_mux2_1
X_4223_ net1192 net1045 _2564_ VPWR VGND sg13g2_nor2b_1
X_4154_ net1225 net1200 _2504_ VPWR VGND sg13g2_nor2b_1
XFILLER_29_919 VPWR VGND sg13g2_decap_4
X_4085_ VPWR _2444_ net326 VGND sg13g2_inv_1
XFILLER_37_985 VPWR VGND sg13g2_decap_8
XFILLER_36_451 VPWR VGND sg13g2_fill_1
X_6066__214 VPWR VGND net214 sg13g2_tiehi
XFILLER_23_101 VPWR VGND sg13g2_decap_8
XFILLER_24_624 VPWR VGND sg13g2_fill_2
X_4987_ VGND VPWR _0614_ _0693_ _0694_ net1140 sg13g2_a21oi_1
X_3938_ net1293 VPWR _2316_ VGND net928 _2315_ sg13g2_o21ai_1
X_3869_ _2253_ net954 _2227_ _2254_ VPWR VGND sg13g2_a21o_1
X_5608_ _1258_ VPWR _1259_ VGND _1254_ _1257_ sg13g2_o21ai_1
X_5539_ _1195_ net1078 _1148_ _1196_ VPWR VGND sg13g2_a21o_1
Xfanout1329 net1331 net1329 VPWR VGND sg13g2_buf_8
Xfanout1318 net1319 net1318 VPWR VGND sg13g2_buf_8
Xfanout1307 net1310 net1307 VPWR VGND sg13g2_buf_8
XFILLER_47_738 VPWR VGND sg13g2_decap_8
XFILLER_4_1019 VPWR VGND sg13g2_decap_8
XFILLER_19_429 VPWR VGND sg13g2_decap_4
XFILLER_36_64 VPWR VGND sg13g2_decap_4
XFILLER_27_440 VPWR VGND sg13g2_decap_8
XFILLER_43_933 VPWR VGND sg13g2_decap_8
XFILLER_27_484 VPWR VGND sg13g2_decap_4
XFILLER_42_498 VPWR VGND sg13g2_decap_4
XFILLER_30_616 VPWR VGND sg13g2_decap_4
XFILLER_11_874 VPWR VGND sg13g2_decap_8
XFILLER_10_384 VPWR VGND sg13g2_decap_8
XFILLER_6_377 VPWR VGND sg13g2_fill_1
XFILLER_6_355 VPWR VGND sg13g2_decap_4
XFILLER_35_7 VPWR VGND sg13g2_fill_1
XFILLER_2_594 VPWR VGND sg13g2_decap_8
XFILLER_18_440 VPWR VGND sg13g2_decap_8
XFILLER_18_451 VPWR VGND sg13g2_fill_1
XFILLER_46_782 VPWR VGND sg13g2_decap_8
X_5890_ net1016 net1059 _1508_ VPWR VGND sg13g2_nor2b_1
X_4910_ s0.data_out\[16\]\[4\] s0.data_out\[15\]\[4\] net1141 _0627_ VPWR VGND sg13g2_mux2_1
XFILLER_33_421 VPWR VGND sg13g2_decap_4
X_4841_ VPWR _0066_ _0562_ VGND sg13g2_inv_1
XFILLER_34_977 VPWR VGND sg13g2_decap_8
X_5983__32 VPWR VGND net32 sg13g2_tiehi
X_4772_ s0.data_out\[17\]\[7\] s0.data_out\[16\]\[7\] net1151 _0501_ VPWR VGND sg13g2_mux2_1
X_3723_ _2076_ VPWR _2120_ VGND net932 _2119_ sg13g2_o21ai_1
X_3654_ VGND VPWR _2443_ _2054_ _0224_ _2060_ sg13g2_a21oi_1
X_3585_ net974 net1046 _1995_ VPWR VGND sg13g2_nor2b_1
XFILLER_0_509 VPWR VGND sg13g2_decap_8
X_5324_ _1002_ VPWR _1003_ VGND net1092 _0996_ sg13g2_o21ai_1
X_5255_ _0937_ s0.data_out\[12\]\[7\] net1121 VPWR VGND sg13g2_nand2b_1
X_4206_ net1196 s0.data_out\[20\]\[5\] _2549_ VPWR VGND sg13g2_and2_1
X_5186_ net1338 net298 _0096_ VPWR VGND sg13g2_and2_1
X_4137_ _2495_ VPWR net2 VGND _2482_ net913 sg13g2_o21ai_1
XFILLER_44_708 VPWR VGND sg13g2_decap_8
X_4068_ net1281 _2399_ _2400_ _2429_ VPWR VGND sg13g2_nor3_1
XFILLER_37_782 VPWR VGND sg13g2_decap_8
XFILLER_25_999 VPWR VGND sg13g2_decap_8
XFILLER_12_638 VPWR VGND sg13g2_fill_1
XFILLER_4_837 VPWR VGND sg13g2_decap_8
Xfanout1104 s0.shift_out\[12\][0] net1104 VPWR VGND sg13g2_buf_2
Xfanout1115 net1116 net1115 VPWR VGND sg13g2_buf_1
Xfanout1126 net1129 net1126 VPWR VGND sg13g2_buf_1
Xfanout1137 net1140 net1137 VPWR VGND sg13g2_buf_1
XFILLER_47_30 VPWR VGND sg13g2_fill_1
Xfanout1159 net1162 net1159 VPWR VGND sg13g2_buf_1
Xfanout1148 net1150 net1148 VPWR VGND sg13g2_buf_8
XFILLER_47_96 VPWR VGND sg13g2_fill_1
XFILLER_35_719 VPWR VGND sg13g2_fill_1
XFILLER_28_782 VPWR VGND sg13g2_decap_4
XFILLER_15_421 VPWR VGND sg13g2_fill_2
XFILLER_30_435 VPWR VGND sg13g2_decap_8
X_5980__35 VPWR VGND net35 sg13g2_tiehi
XFILLER_11_660 VPWR VGND sg13g2_fill_2
XFILLER_8_79 VPWR VGND sg13g2_fill_1
XFILLER_8_68 VPWR VGND sg13g2_decap_8
XFILLER_7_686 VPWR VGND sg13g2_decap_4
X_3370_ _1802_ VPWR _1803_ VGND net1264 _1784_ sg13g2_o21ai_1
X_5040_ _0680_ VPWR _0745_ VGND _2464_ _0744_ sg13g2_o21ai_1
XFILLER_33_4 VPWR VGND sg13g2_fill_2
XFILLER_19_760 VPWR VGND sg13g2_decap_8
X_5942_ _1556_ net1020 net544 VPWR VGND sg13g2_nand2_1
XFILLER_18_281 VPWR VGND sg13g2_fill_2
X_6063__217 VPWR VGND net217 sg13g2_tiehi
XFILLER_22_914 VPWR VGND sg13g2_fill_2
X_5873_ net1013 net1067 _1493_ VPWR VGND sg13g2_nor2b_1
X_4824_ _0547_ VPWR _0548_ VGND net1317 net476 sg13g2_o21ai_1
X_4755_ s0.data_out\[17\]\[0\] s0.data_out\[16\]\[0\] net1151 _0484_ VPWR VGND sg13g2_mux2_1
X_3706_ net964 net1050 _2105_ VPWR VGND sg13g2_nor2b_1
X_4686_ net1144 s0.data_out\[16\]\[0\] _0423_ VPWR VGND sg13g2_and2_1
X_3637_ _2036_ VPWR _2046_ VGND _2041_ _2043_ sg13g2_o21ai_1
X_3568_ _1980_ _2471_ _1979_ VPWR VGND sg13g2_nand2_1
X_5307_ net1251 _0986_ _0988_ VPWR VGND sg13g2_nor2_1
X_3499_ VGND VPWR net984 _1919_ _1920_ _1865_ sg13g2_a21oi_1
X_5238_ VPWR _0103_ _0922_ VGND sg13g2_inv_1
XFILLER_25_1020 VPWR VGND sg13g2_decap_8
X_5169_ _0862_ net1121 net599 VPWR VGND sg13g2_nand2_1
XFILLER_40_711 VPWR VGND sg13g2_fill_1
XFILLER_25_763 VPWR VGND sg13g2_fill_1
XFILLER_12_424 VPWR VGND sg13g2_fill_1
XFILLER_12_435 VPWR VGND sg13g2_decap_8
XFILLER_12_446 VPWR VGND sg13g2_fill_1
XFILLER_24_295 VPWR VGND sg13g2_decap_4
XFILLER_9_929 VPWR VGND sg13g2_decap_8
XFILLER_12_479 VPWR VGND sg13g2_fill_2
XFILLER_32_1024 VPWR VGND sg13g2_decap_4
XFILLER_0_873 VPWR VGND sg13g2_decap_8
XFILLER_48_822 VPWR VGND sg13g2_decap_8
Xhold6 s0.genblk1\[12\].modules.bubble VPWR VGND net302 sg13g2_dlygate4sd3_1
XFILLER_48_899 VPWR VGND sg13g2_decap_8
XFILLER_16_752 VPWR VGND sg13g2_fill_1
XFILLER_28_590 VPWR VGND sg13g2_decap_8
XFILLER_30_254 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_10_clk clknet_3_2__leaf_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
X_4540_ VGND VPWR _0293_ net1208 net305 sg13g2_or2_1
XFILLER_7_472 VPWR VGND sg13g2_decap_4
X_4471_ VPWR _0032_ _2789_ VGND sg13g2_inv_1
X_6210_ net234 VGND VPWR _0260_ s0.was_valid_out\[0\][0] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_3422_ s0.data_out\[4\]\[3\] s0.data_out\[5\]\[3\] net997 _1848_ VPWR VGND sg13g2_mux2_1
X_6141_ net133 VGND VPWR _0191_ s0.data_out\[6\]\[1\] clknet_leaf_23_clk sg13g2_dfrbpq_2
Xfanout919 _2466_ net919 VPWR VGND sg13g2_buf_8
X_3353_ _1785_ VPWR _1786_ VGND _1779_ _1780_ sg13g2_o21ai_1
X_6072_ net207 VGND VPWR _0122_ s0.valid_out\[11\][0] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_3284_ VGND VPWR _1724_ net537 net1324 sg13g2_or2_1
XFILLER_38_321 VPWR VGND sg13g2_decap_4
X_5023_ _0727_ VPWR _0728_ VGND _0720_ _0721_ sg13g2_o21ai_1
XFILLER_38_376 VPWR VGND sg13g2_fill_1
X_5925_ VGND VPWR net1023 _1538_ _1539_ _1485_ sg13g2_a21oi_1
X_5856_ _1478_ net918 _1477_ VPWR VGND sg13g2_nand2_1
X_4807_ net1319 VPWR _0534_ VGND _0531_ _0533_ sg13g2_o21ai_1
X_5787_ VPWR _0161_ net566 VGND sg13g2_inv_1
XFILLER_21_276 VPWR VGND sg13g2_fill_2
X_4738_ _0468_ VPWR _0469_ VGND _0464_ _0467_ sg13g2_o21ai_1
X_4669_ _0298_ _0408_ _0409_ _0410_ VPWR VGND sg13g2_nor3_1
XFILLER_1_648 VPWR VGND sg13g2_decap_8
XFILLER_0_158 VPWR VGND sg13g2_decap_8
XFILLER_44_313 VPWR VGND sg13g2_fill_1
XFILLER_45_858 VPWR VGND sg13g2_decap_8
XFILLER_40_530 VPWR VGND sg13g2_decap_8
XFILLER_13_733 VPWR VGND sg13g2_decap_8
XFILLER_25_571 VPWR VGND sg13g2_fill_1
XFILLER_12_243 VPWR VGND sg13g2_decap_8
XFILLER_12_254 VPWR VGND sg13g2_fill_2
XFILLER_40_585 VPWR VGND sg13g2_fill_2
XFILLER_8_269 VPWR VGND sg13g2_fill_1
XFILLER_8_258 VPWR VGND sg13g2_decap_8
XFILLER_5_965 VPWR VGND sg13g2_decap_8
XFILLER_4_431 VPWR VGND sg13g2_decap_8
XFILLER_0_670 VPWR VGND sg13g2_decap_8
XFILLER_48_696 VPWR VGND sg13g2_decap_8
XFILLER_35_324 VPWR VGND sg13g2_fill_2
X_3971_ VGND VPWR _2345_ net495 net1299 sg13g2_or2_1
XFILLER_23_508 VPWR VGND sg13g2_fill_1
X_5710_ VGND VPWR net1223 _2474_ _0150_ _1347_ sg13g2_a21oi_1
X_5641_ VPWR _0141_ net522 VGND sg13g2_inv_1
XFILLER_31_596 VPWR VGND sg13g2_fill_1
X_5572_ VGND VPWR _1224_ _1227_ _0131_ _1228_ sg13g2_a21oi_1
X_4523_ _0275_ net1172 _2785_ _0276_ VPWR VGND sg13g2_a21o_1
Xhold225 s0.data_out\[10\]\[6\] VPWR VGND net521 sg13g2_dlygate4sd3_1
Xhold203 _0324_ VPWR VGND net499 sg13g2_dlygate4sd3_1
Xhold214 _2088_ VPWR VGND net510 sg13g2_dlygate4sd3_1
Xhold247 _1406_ VPWR VGND net543 sg13g2_dlygate4sd3_1
Xhold269 s0.data_out\[9\]\[7\] VPWR VGND net565 sg13g2_dlygate4sd3_1
Xhold236 _1294_ VPWR VGND net532 sg13g2_dlygate4sd3_1
X_4454_ _2774_ VPWR _2775_ VGND _2770_ _2773_ sg13g2_o21ai_1
Xhold258 s0.data_out\[15\]\[7\] VPWR VGND net554 sg13g2_dlygate4sd3_1
X_4385_ _2713_ net1188 net551 VPWR VGND sg13g2_nand2_1
X_3405_ VPWR _0202_ _1833_ VGND sg13g2_inv_1
X_6124_ net152 VGND VPWR _0174_ s0.shift_out\[8\][0] clknet_leaf_16_clk sg13g2_dfrbpq_2
X_3336_ s0.data_out\[6\]\[2\] s0.data_out\[5\]\[2\] net999 _1769_ VPWR VGND sg13g2_mux2_1
X_6055_ net226 VGND VPWR _0105_ s0.data_out\[13\]\[6\] clknet_leaf_27_clk sg13g2_dfrbpq_2
X_3267_ VGND VPWR _1704_ _1707_ _1710_ _1709_ sg13g2_a21oi_1
X_5006_ _0710_ _0666_ net1271 _0711_ VPWR VGND sg13g2_a21o_1
X_3198_ VGND VPWR _1552_ _1643_ _1644_ net1018 sg13g2_a21oi_1
XFILLER_38_173 VPWR VGND sg13g2_fill_1
XFILLER_38_195 VPWR VGND sg13g2_decap_8
XFILLER_27_858 VPWR VGND sg13g2_decap_8
XFILLER_27_869 VPWR VGND sg13g2_fill_2
XFILLER_14_508 VPWR VGND sg13g2_fill_2
XFILLER_41_338 VPWR VGND sg13g2_decap_8
XFILLER_41_327 VPWR VGND sg13g2_fill_2
X_5908_ VGND VPWR _1524_ net587 net1330 sg13g2_or2_1
X_5839_ _1454_ VPWR _1465_ VGND _1458_ _1460_ sg13g2_o21ai_1
XFILLER_10_725 VPWR VGND sg13g2_decap_8
XFILLER_6_718 VPWR VGND sg13g2_decap_8
XFILLER_5_206 VPWR VGND sg13g2_decap_8
XFILLER_5_239 VPWR VGND sg13g2_fill_2
XFILLER_2_924 VPWR VGND sg13g2_decap_8
XFILLER_7_1006 VPWR VGND sg13g2_decap_8
XFILLER_29_140 VPWR VGND sg13g2_fill_1
XFILLER_29_151 VPWR VGND sg13g2_decap_8
XFILLER_29_195 VPWR VGND sg13g2_decap_8
XFILLER_32_349 VPWR VGND sg13g2_fill_1
XFILLER_41_883 VPWR VGND sg13g2_decap_4
XFILLER_9_523 VPWR VGND sg13g2_fill_1
XFILLER_13_585 VPWR VGND sg13g2_fill_1
XFILLER_40_393 VPWR VGND sg13g2_decap_8
XFILLER_40_382 VPWR VGND sg13g2_fill_1
XFILLER_45_1012 VPWR VGND sg13g2_decap_8
X_4170_ net1206 s0.data_out\[20\]\[0\] _2518_ VPWR VGND sg13g2_nor2_1
X_3121_ _1568_ _1574_ _1551_ _1578_ VPWR VGND _1577_ sg13g2_nand4_1
XFILLER_49_961 VPWR VGND sg13g2_decap_8
XFILLER_48_471 VPWR VGND sg13g2_decap_8
XFILLER_36_666 VPWR VGND sg13g2_fill_2
XFILLER_35_165 VPWR VGND sg13g2_fill_2
XFILLER_35_154 VPWR VGND sg13g2_fill_2
XFILLER_17_880 VPWR VGND sg13g2_fill_2
X_3954_ net952 VPWR _2330_ VGND _2328_ _2329_ sg13g2_o21ai_1
XFILLER_32_861 VPWR VGND sg13g2_decap_8
X_3885_ VGND VPWR net953 _2269_ _2270_ _2214_ sg13g2_a21oi_1
X_5624_ _1272_ VPWR _1273_ VGND net1344 net429 sg13g2_o21ai_1
X_6105__172 VPWR VGND net172 sg13g2_tiehi
X_5555_ _1211_ net1081 _1155_ _1212_ VPWR VGND sg13g2_a21o_1
X_4506_ _2822_ net1262 _2821_ VPWR VGND sg13g2_nand2_1
X_5486_ net1079 net1062 _1148_ VPWR VGND sg13g2_nor2b_1
XFILLER_6_90 VPWR VGND sg13g2_fill_2
X_4437_ _2756_ _2759_ net1302 _2760_ VPWR VGND sg13g2_nand3_1
X_4368_ _2696_ net1193 _2695_ VPWR VGND sg13g2_nand2b_1
X_6107_ net170 VGND VPWR _0157_ s0.data_out\[9\]\[3\] clknet_leaf_22_clk sg13g2_dfrbpq_2
X_3319_ _1754_ net538 net1009 VPWR VGND sg13g2_nand2b_1
X_4299_ net1178 s0.data_out\[19\]\[0\] _2635_ VPWR VGND sg13g2_and2_1
X_6038_ net244 VGND VPWR _0088_ s0.data_out\[14\]\[1\] clknet_leaf_29_clk sg13g2_dfrbpq_2
X_6112__165 VPWR VGND net165 sg13g2_tiehi
XFILLER_25_11 VPWR VGND sg13g2_decap_8
XFILLER_23_861 VPWR VGND sg13g2_decap_4
XFILLER_10_533 VPWR VGND sg13g2_decap_8
XFILLER_2_721 VPWR VGND sg13g2_decap_8
XFILLER_2_798 VPWR VGND sg13g2_decap_8
XFILLER_37_408 VPWR VGND sg13g2_fill_1
XFILLER_18_611 VPWR VGND sg13g2_decap_4
XFILLER_17_110 VPWR VGND sg13g2_decap_8
XFILLER_46_964 VPWR VGND sg13g2_decap_8
XFILLER_17_143 VPWR VGND sg13g2_decap_4
XFILLER_17_154 VPWR VGND sg13g2_decap_8
XFILLER_33_603 VPWR VGND sg13g2_fill_1
XFILLER_45_474 VPWR VGND sg13g2_decap_8
XFILLER_33_614 VPWR VGND sg13g2_fill_1
XFILLER_33_625 VPWR VGND sg13g2_fill_1
XFILLER_33_647 VPWR VGND sg13g2_fill_1
XFILLER_9_342 VPWR VGND sg13g2_fill_2
X_3670_ _2073_ VPWR _2074_ VGND net1307 net421 sg13g2_o21ai_1
X_6059__222 VPWR VGND net222 sg13g2_tiehi
X_5340_ VGND VPWR net1088 s0.data_out\[11\]\[1\] _1016_ _1015_ sg13g2_a21oi_1
XFILLER_5_581 VPWR VGND sg13g2_decap_8
X_5271_ _0896_ _0951_ net1279 _0952_ VPWR VGND sg13g2_nand3_1
X_4222_ net1192 s0.data_out\[20\]\[7\] _2563_ VPWR VGND sg13g2_and2_1
X_4153_ net1204 VPWR _2503_ VGND net1225 net1195 sg13g2_o21ai_1
X_4084_ VPWR _2443_ net319 VGND sg13g2_inv_1
XFILLER_37_964 VPWR VGND sg13g2_decap_8
XFILLER_36_463 VPWR VGND sg13g2_fill_2
X_4986_ _0693_ s0.data_out\[14\]\[6\] net1142 VPWR VGND sg13g2_nand2b_1
XFILLER_24_647 VPWR VGND sg13g2_fill_2
XFILLER_23_179 VPWR VGND sg13g2_decap_4
X_3937_ VGND VPWR net941 net348 _2315_ _2314_ sg13g2_a21oi_1
X_3868_ s0.data_out\[2\]\[7\] s0.data_out\[1\]\[7\] net957 _2253_ VPWR VGND sg13g2_mux2_1
XFILLER_20_853 VPWR VGND sg13g2_decap_8
X_5607_ VGND VPWR _1258_ net506 net1344 sg13g2_or2_1
X_3799_ _2190_ net458 net965 VPWR VGND sg13g2_nand2b_1
XFILLER_11_57 VPWR VGND sg13g2_fill_2
X_5538_ s0.data_out\[11\]\[3\] s0.data_out\[10\]\[3\] net1084 _1195_ VPWR VGND sg13g2_mux2_1
X_5469_ VGND VPWR _1067_ _1132_ _1133_ net1090 sg13g2_a21oi_1
Xfanout1319 net1323 net1319 VPWR VGND sg13g2_buf_8
Xfanout1308 net1310 net1308 VPWR VGND sg13g2_buf_1
XFILLER_47_717 VPWR VGND sg13g2_decap_8
XFILLER_46_249 VPWR VGND sg13g2_fill_2
XFILLER_43_912 VPWR VGND sg13g2_decap_8
XFILLER_28_986 VPWR VGND sg13g2_decap_8
XFILLER_43_989 VPWR VGND sg13g2_decap_8
XFILLER_11_831 VPWR VGND sg13g2_fill_2
XFILLER_7_824 VPWR VGND sg13g2_fill_1
XFILLER_11_886 VPWR VGND sg13g2_decap_4
XFILLER_6_334 VPWR VGND sg13g2_decap_8
XFILLER_38_739 VPWR VGND sg13g2_decap_8
XFILLER_19_920 VPWR VGND sg13g2_decap_8
XFILLER_46_761 VPWR VGND sg13g2_decap_8
X_4840_ _0561_ VPWR _0562_ VGND _0557_ _0560_ sg13g2_o21ai_1
XFILLER_34_956 VPWR VGND sg13g2_decap_8
XFILLER_33_466 VPWR VGND sg13g2_fill_2
X_4771_ _0500_ net1152 net591 VPWR VGND sg13g2_nand2_1
XFILLER_20_116 VPWR VGND sg13g2_fill_1
XFILLER_33_499 VPWR VGND sg13g2_fill_2
XFILLER_9_150 VPWR VGND sg13g2_decap_4
X_3722_ VGND VPWR net959 _2118_ _2119_ _2078_ sg13g2_a21oi_1
X_3653_ net1309 VPWR _2060_ VGND _2057_ _2059_ sg13g2_o21ai_1
X_3584_ VGND VPWR _1903_ _1993_ _1994_ net983 sg13g2_a21oi_1
X_5323_ net938 VPWR _1002_ VGND s0.was_valid_out\[11\][0] net1110 sg13g2_o21ai_1
X_5254_ VPWR _0105_ _0936_ VGND sg13g2_inv_1
X_5185_ VGND VPWR _0872_ _0876_ _0095_ _0877_ sg13g2_a21oi_1
X_4205_ _0007_ _2544_ _2548_ _2477_ net1217 VPWR VGND sg13g2_a22oi_1
X_4136_ _2495_ net1281 net913 VPWR VGND sg13g2_nand2_1
XFILLER_29_706 VPWR VGND sg13g2_fill_2
XFILLER_3_1020 VPWR VGND sg13g2_decap_8
XFILLER_28_238 VPWR VGND sg13g2_decap_8
XFILLER_25_901 VPWR VGND sg13g2_fill_2
X_4067_ net1274 VPWR _2428_ VGND _2402_ _2403_ sg13g2_o21ai_1
XFILLER_40_959 VPWR VGND sg13g2_decap_8
X_4969_ VPWR _0078_ _0678_ VGND sg13g2_inv_1
XFILLER_20_683 VPWR VGND sg13g2_decap_8
XFILLER_4_816 VPWR VGND sg13g2_decap_8
XFILLER_22_89 VPWR VGND sg13g2_fill_1
XFILLER_3_315 VPWR VGND sg13g2_fill_1
Xfanout1116 net1118 net1116 VPWR VGND sg13g2_buf_8
Xfanout1127 net1128 net1127 VPWR VGND sg13g2_buf_8
Xfanout1138 net1139 net1138 VPWR VGND sg13g2_buf_8
Xfanout1105 net1106 net1105 VPWR VGND sg13g2_buf_8
Xfanout1149 net1150 net1149 VPWR VGND sg13g2_buf_8
XFILLER_19_238 VPWR VGND sg13g2_decap_8
X_6049__232 VPWR VGND net232 sg13g2_tiehi
XFILLER_15_433 VPWR VGND sg13g2_decap_8
XFILLER_16_945 VPWR VGND sg13g2_fill_2
XFILLER_27_282 VPWR VGND sg13g2_decap_8
XFILLER_42_263 VPWR VGND sg13g2_fill_1
XFILLER_15_477 VPWR VGND sg13g2_fill_1
X_6056__225 VPWR VGND net225 sg13g2_tiehi
XFILLER_26_4 VPWR VGND sg13g2_decap_8
X_5941_ VGND VPWR net1025 _1554_ _1555_ _1527_ sg13g2_a21oi_1
XFILLER_18_293 VPWR VGND sg13g2_decap_8
X_5872_ VGND VPWR _1414_ _1491_ _1492_ net1024 sg13g2_a21oi_1
XFILLER_33_241 VPWR VGND sg13g2_decap_4
XFILLER_34_775 VPWR VGND sg13g2_fill_2
X_4823_ _0543_ _0546_ net1317 _0547_ VPWR VGND sg13g2_nand3_1
XFILLER_21_425 VPWR VGND sg13g2_decap_4
XFILLER_22_959 VPWR VGND sg13g2_fill_1
X_4754_ VGND VPWR net1160 _0482_ _0483_ _0429_ sg13g2_a21oi_1
XFILLER_21_458 VPWR VGND sg13g2_decap_4
X_3705_ VGND VPWR _2024_ _2103_ _2104_ net973 sg13g2_a21oi_1
XFILLER_30_981 VPWR VGND sg13g2_decap_8
X_4685_ _0422_ net924 _0421_ VPWR VGND sg13g2_nand2_1
X_3636_ _2031_ _2044_ _2019_ _2045_ VPWR VGND sg13g2_nand3_1
X_3567_ s0.data_out\[3\]\[5\] s0.data_out\[4\]\[5\] net988 _1979_ VPWR VGND sg13g2_mux2_1
X_5306_ _0987_ net1251 _0986_ VPWR VGND sg13g2_nand2_1
X_3498_ s0.data_out\[5\]\[5\] s0.data_out\[4\]\[5\] net989 _1919_ VPWR VGND sg13g2_mux2_1
XFILLER_0_329 VPWR VGND sg13g2_decap_8
X_5237_ _0921_ VPWR _0922_ VGND net1334 net430 sg13g2_o21ai_1
X_5168_ _0861_ net1256 _0860_ VPWR VGND sg13g2_nand2_1
X_4119_ VPWR _2478_ net366 VGND sg13g2_inv_1
X_5099_ _0793_ _0796_ net1321 _0797_ VPWR VGND sg13g2_nand3_1
XFILLER_44_517 VPWR VGND sg13g2_fill_2
XFILLER_25_775 VPWR VGND sg13g2_fill_2
XFILLER_40_745 VPWR VGND sg13g2_fill_2
XFILLER_33_33 VPWR VGND sg13g2_fill_2
XFILLER_40_778 VPWR VGND sg13g2_decap_4
XFILLER_32_1003 VPWR VGND sg13g2_decap_8
XFILLER_33_88 VPWR VGND sg13g2_fill_1
XFILLER_4_613 VPWR VGND sg13g2_decap_8
XFILLER_4_679 VPWR VGND sg13g2_decap_8
XFILLER_48_801 VPWR VGND sg13g2_decap_8
XFILLER_0_852 VPWR VGND sg13g2_decap_8
Xhold7 s0.genblk1\[14\].modules.bubble VPWR VGND net303 sg13g2_dlygate4sd3_1
XFILLER_48_878 VPWR VGND sg13g2_decap_8
XFILLER_47_377 VPWR VGND sg13g2_fill_2
XFILLER_15_274 VPWR VGND sg13g2_decap_4
XFILLER_12_992 VPWR VGND sg13g2_decap_8
XFILLER_8_985 VPWR VGND sg13g2_decap_8
X_4470_ _2788_ VPWR _2789_ VGND _2784_ _2787_ sg13g2_o21ai_1
X_3421_ VPWR _0204_ _1847_ VGND sg13g2_inv_1
X_6140_ net134 VGND VPWR _0190_ s0.data_out\[6\]\[0\] clknet_leaf_23_clk sg13g2_dfrbpq_2
X_3352_ _1785_ _1784_ net1264 _1771_ net1271 VPWR VGND sg13g2_a22oi_1
X_6071_ net209 VGND VPWR _0121_ s0.was_valid_out\[11\][0] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_3283_ net1324 VPWR _1723_ VGND net916 _1722_ sg13g2_o21ai_1
X_5022_ VGND VPWR net1264 _0726_ _0727_ _0722_ sg13g2_a21oi_1
XFILLER_17_0 VPWR VGND sg13g2_fill_2
XFILLER_0_92 VPWR VGND sg13g2_fill_1
X_5924_ _1537_ net1013 _1486_ _1538_ VPWR VGND sg13g2_a21o_1
X_5855_ s0.data_out\[7\]\[0\] s0.data_out\[8\]\[0\] net1031 _1477_ VPWR VGND sg13g2_mux2_1
X_4806_ _0533_ _0530_ _0532_ VPWR VGND sg13g2_nand2_1
XFILLER_21_222 VPWR VGND sg13g2_fill_1
XFILLER_21_233 VPWR VGND sg13g2_fill_2
XFILLER_22_778 VPWR VGND sg13g2_decap_4
X_5786_ _1412_ VPWR _1413_ VGND _1408_ _1411_ sg13g2_o21ai_1
X_4737_ VGND VPWR _0468_ net572 net1304 sg13g2_or2_1
X_4668_ _0389_ _0391_ _0409_ VPWR VGND sg13g2_nor2b_1
X_3619_ _2028_ _2027_ net1241 _2023_ net1233 VPWR VGND sg13g2_a22oi_1
X_4599_ net1303 VPWR _0343_ VGND _2461_ _0342_ sg13g2_o21ai_1
XFILLER_0_104 VPWR VGND sg13g2_decap_4
XFILLER_1_627 VPWR VGND sg13g2_decap_8
XFILLER_45_837 VPWR VGND sg13g2_decap_8
XFILLER_29_377 VPWR VGND sg13g2_fill_1
XFILLER_29_388 VPWR VGND sg13g2_decap_8
XFILLER_44_87 VPWR VGND sg13g2_decap_4
XFILLER_44_76 VPWR VGND sg13g2_fill_1
XFILLER_25_594 VPWR VGND sg13g2_fill_1
XFILLER_9_716 VPWR VGND sg13g2_decap_8
XFILLER_40_564 VPWR VGND sg13g2_fill_2
XFILLER_8_237 VPWR VGND sg13g2_decap_8
XFILLER_8_226 VPWR VGND sg13g2_fill_1
XFILLER_5_944 VPWR VGND sg13g2_decap_8
XFILLER_4_465 VPWR VGND sg13g2_fill_2
X_6053__228 VPWR VGND net228 sg13g2_tiehi
XFILLER_48_675 VPWR VGND sg13g2_decap_8
XFILLER_36_859 VPWR VGND sg13g2_fill_2
XFILLER_36_848 VPWR VGND sg13g2_decap_8
X_3970_ net1295 VPWR _2344_ VGND net929 _2343_ sg13g2_o21ai_1
XFILLER_44_892 VPWR VGND sg13g2_decap_8
XFILLER_31_520 VPWR VGND sg13g2_decap_4
XFILLER_43_391 VPWR VGND sg13g2_decap_4
X_5640_ _1286_ VPWR _1287_ VGND _1282_ _1285_ sg13g2_o21ai_1
X_5571_ VGND VPWR _1228_ net1210 net316 sg13g2_or2_1
X_4522_ s0.data_out\[19\]\[5\] s0.data_out\[18\]\[5\] net1176 _0275_ VPWR VGND sg13g2_mux2_1
Xhold215 s0.data_out\[4\]\[6\] VPWR VGND net511 sg13g2_dlygate4sd3_1
Xhold226 _1287_ VPWR VGND net522 sg13g2_dlygate4sd3_1
XFILLER_8_793 VPWR VGND sg13g2_fill_1
X_4453_ VGND VPWR _2774_ net567 net1287 sg13g2_or2_1
Xhold204 s0.valid_out\[11\][0] VPWR VGND net500 sg13g2_dlygate4sd3_1
Xhold248 s0.data_out\[7\]\[6\] VPWR VGND net544 sg13g2_dlygate4sd3_1
Xhold259 _0706_ VPWR VGND net555 sg13g2_dlygate4sd3_1
X_3404_ _1832_ VPWR _1833_ VGND net1311 net432 sg13g2_o21ai_1
Xhold237 s0.data_out\[4\]\[2\] VPWR VGND net533 sg13g2_dlygate4sd3_1
X_4384_ VGND VPWR net1197 _2711_ _2712_ _2683_ sg13g2_a21oi_1
X_6123_ net153 VGND VPWR _0173_ s0.data_out\[8\]\[7\] clknet_leaf_18_clk sg13g2_dfrbpq_2
X_3335_ _1768_ net997 net581 VPWR VGND sg13g2_nand2_1
X_3266_ _1708_ VPWR _1709_ VGND net995 _1702_ sg13g2_o21ai_1
X_6054_ net227 VGND VPWR _0104_ s0.data_out\[13\]\[5\] clknet_leaf_28_clk sg13g2_dfrbpq_2
X_5005_ _0710_ net1138 _0709_ VPWR VGND sg13g2_nand2b_1
XFILLER_22_1013 VPWR VGND sg13g2_decap_8
X_3197_ _1643_ s0.data_out\[6\]\[7\] net1021 VPWR VGND sg13g2_nand2b_1
XFILLER_39_664 VPWR VGND sg13g2_fill_1
XFILLER_38_185 VPWR VGND sg13g2_decap_4
XFILLER_26_347 VPWR VGND sg13g2_fill_1
X_5907_ net1330 VPWR _1523_ VGND net918 _1522_ sg13g2_o21ai_1
XFILLER_34_380 VPWR VGND sg13g2_fill_2
X_5838_ _1449_ _1459_ _1435_ _1464_ VPWR VGND _1463_ sg13g2_nand4_1
XFILLER_14_68 VPWR VGND sg13g2_fill_2
X_5769_ _1394_ _1397_ net1342 _1398_ VPWR VGND sg13g2_nand3_1
XFILLER_2_903 VPWR VGND sg13g2_decap_8
XFILLER_39_65 VPWR VGND sg13g2_fill_2
XFILLER_18_815 VPWR VGND sg13g2_fill_1
XFILLER_18_848 VPWR VGND sg13g2_fill_1
XFILLER_17_358 VPWR VGND sg13g2_fill_2
XFILLER_33_807 VPWR VGND sg13g2_fill_1
XFILLER_44_166 VPWR VGND sg13g2_fill_2
XFILLER_26_892 VPWR VGND sg13g2_decap_8
XFILLER_25_380 VPWR VGND sg13g2_decap_4
XFILLER_9_502 VPWR VGND sg13g2_fill_2
X_3120_ _1563_ _1575_ _1576_ _1577_ VPWR VGND sg13g2_nor3_1
XFILLER_49_940 VPWR VGND sg13g2_decap_8
XFILLER_1_991 VPWR VGND sg13g2_decap_8
XFILLER_48_450 VPWR VGND sg13g2_decap_8
XFILLER_35_133 VPWR VGND sg13g2_decap_4
X_3953_ net943 net1053 _2329_ VPWR VGND sg13g2_nor2b_1
X_3884_ s0.data_out\[2\]\[5\] s0.data_out\[1\]\[5\] net957 _2269_ VPWR VGND sg13g2_mux2_1
X_5623_ _1268_ _1271_ net1344 _1272_ VPWR VGND sg13g2_nand3_1
X_5554_ s0.data_out\[11\]\[4\] s0.data_out\[10\]\[4\] net1085 _1211_ VPWR VGND sg13g2_mux2_1
X_4505_ VGND VPWR net1181 _2820_ _2821_ _2770_ sg13g2_a21oi_1
X_5485_ VGND VPWR _1077_ _1146_ _1147_ net1090 sg13g2_a21oi_1
X_4436_ net1181 VPWR _2759_ VGND _2757_ _2758_ sg13g2_o21ai_1
X_4367_ VGND VPWR net1178 _2694_ _2695_ _2643_ sg13g2_a21oi_1
X_3318_ VPWR _0195_ _1753_ VGND sg13g2_inv_1
X_6106_ net171 VGND VPWR _0156_ s0.data_out\[9\]\[2\] clknet_leaf_22_clk sg13g2_dfrbpq_2
X_4298_ _2634_ net931 _2633_ VPWR VGND sg13g2_nand2_1
X_3249_ VGND VPWR _1694_ _1686_ net1238 sg13g2_or2_1
X_6037_ net245 VGND VPWR _0087_ s0.data_out\[14\]\[0\] clknet_leaf_30_clk sg13g2_dfrbpq_2
XFILLER_26_100 VPWR VGND sg13g2_decap_4
XFILLER_15_818 VPWR VGND sg13g2_decap_4
XFILLER_42_626 VPWR VGND sg13g2_fill_2
XFILLER_41_114 VPWR VGND sg13g2_decap_4
XFILLER_25_34 VPWR VGND sg13g2_fill_1
XFILLER_25_45 VPWR VGND sg13g2_decap_4
XFILLER_41_169 VPWR VGND sg13g2_decap_8
XFILLER_41_158 VPWR VGND sg13g2_fill_1
XFILLER_2_700 VPWR VGND sg13g2_decap_8
XFILLER_49_203 VPWR VGND sg13g2_decap_8
XFILLER_2_777 VPWR VGND sg13g2_decap_8
XFILLER_46_943 VPWR VGND sg13g2_decap_8
XFILLER_45_420 VPWR VGND sg13g2_fill_2
XFILLER_32_125 VPWR VGND sg13g2_decap_8
XFILLER_13_361 VPWR VGND sg13g2_decap_4
XFILLER_14_862 VPWR VGND sg13g2_fill_2
XFILLER_14_873 VPWR VGND sg13g2_fill_1
XFILLER_14_884 VPWR VGND sg13g2_decap_8
XFILLER_41_681 VPWR VGND sg13g2_decap_4
XFILLER_13_394 VPWR VGND sg13g2_fill_2
XFILLER_9_398 VPWR VGND sg13g2_fill_1
X_5270_ _0951_ net1116 _0950_ VPWR VGND sg13g2_nand2b_1
X_5998__288 VPWR VGND net288 sg13g2_tiehi
X_4221_ _0009_ _2558_ _2562_ _2473_ net1216 VPWR VGND sg13g2_a22oi_1
X_4152_ net1294 net312 _0000_ VPWR VGND sg13g2_and2_1
X_4083_ VPWR _2442_ net328 VGND sg13g2_inv_1
XFILLER_37_943 VPWR VGND sg13g2_decap_8
XFILLER_37_921 VPWR VGND sg13g2_fill_1
XFILLER_36_442 VPWR VGND sg13g2_decap_8
XFILLER_36_497 VPWR VGND sg13g2_fill_1
X_4985_ VPWR _0080_ _0692_ VGND sg13g2_inv_1
X_3936_ net941 net1061 _2314_ VPWR VGND sg13g2_nor2b_1
X_3867_ _2252_ net956 net495 VPWR VGND sg13g2_nand2_1
XFILLER_20_898 VPWR VGND sg13g2_decap_8
X_3798_ VPWR _0239_ net427 VGND sg13g2_inv_1
X_5606_ net1344 VPWR _1257_ VGND net934 _1256_ sg13g2_o21ai_1
X_5537_ _1185_ _1192_ _1193_ _1194_ VPWR VGND sg13g2_nor3_1
X_5468_ _1132_ net418 net1099 VPWR VGND sg13g2_nand2b_1
Xfanout1309 net1310 net1309 VPWR VGND sg13g2_buf_8
X_4419_ net927 VPWR _2745_ VGND s0.was_valid_out\[18\][0] net1188 sg13g2_o21ai_1
X_5399_ s0.data_out\[12\]\[1\] s0.data_out\[11\]\[1\] net1096 _1068_ VPWR VGND sg13g2_mux2_1
XFILLER_19_409 VPWR VGND sg13g2_decap_4
XFILLER_36_11 VPWR VGND sg13g2_fill_2
XFILLER_28_954 VPWR VGND sg13g2_decap_8
XFILLER_42_401 VPWR VGND sg13g2_fill_2
XFILLER_43_968 VPWR VGND sg13g2_decap_8
XFILLER_14_125 VPWR VGND sg13g2_fill_2
XFILLER_15_648 VPWR VGND sg13g2_decap_8
XFILLER_27_497 VPWR VGND sg13g2_fill_1
XFILLER_11_821 VPWR VGND sg13g2_fill_2
XFILLER_7_803 VPWR VGND sg13g2_decap_4
XFILLER_10_353 VPWR VGND sg13g2_fill_2
XFILLER_2_563 VPWR VGND sg13g2_decap_8
XFILLER_42_1027 VPWR VGND sg13g2_fill_2
XFILLER_38_729 VPWR VGND sg13g2_fill_1
XFILLER_37_228 VPWR VGND sg13g2_decap_8
XFILLER_46_740 VPWR VGND sg13g2_decap_8
XFILLER_45_250 VPWR VGND sg13g2_decap_4
XFILLER_18_475 VPWR VGND sg13g2_fill_2
XFILLER_19_987 VPWR VGND sg13g2_decap_8
XFILLER_34_935 VPWR VGND sg13g2_decap_8
XFILLER_45_283 VPWR VGND sg13g2_decap_8
XFILLER_33_478 VPWR VGND sg13g2_fill_2
X_4770_ VGND VPWR net1161 _0498_ _0499_ _0464_ sg13g2_a21oi_1
X_3721_ _2117_ VPWR _2118_ VGND net968 _2492_ sg13g2_o21ai_1
X_3652_ _2059_ _2056_ _2058_ VPWR VGND sg13g2_nand2_1
X_3583_ _1993_ net515 net988 VPWR VGND sg13g2_nand2b_1
X_6102__176 VPWR VGND net176 sg13g2_tiehi
XFILLER_6_891 VPWR VGND sg13g2_decap_8
X_5322_ VGND VPWR _1001_ net1098 s0.was_valid_out\[11\][0] sg13g2_or2_1
XFILLER_47_0 VPWR VGND sg13g2_decap_8
X_5253_ _0935_ VPWR _0936_ VGND _0931_ _0934_ sg13g2_o21ai_1
X_5184_ VGND VPWR _0877_ net1209 net303 sg13g2_or2_1
X_4204_ net1217 _2547_ _2548_ VPWR VGND sg13g2_nor2_1
XFILLER_3_81 VPWR VGND sg13g2_fill_1
X_4135_ s0.was_valid_out\[21\][0] net1204 _2494_ VPWR VGND sg13g2_nor2_1
X_4066_ _2427_ _2419_ net1246 _2414_ net1254 VPWR VGND sg13g2_a22oi_1
XFILLER_24_434 VPWR VGND sg13g2_decap_8
XFILLER_40_916 VPWR VGND sg13g2_decap_4
XFILLER_40_938 VPWR VGND sg13g2_decap_8
X_4968_ _0677_ VPWR _0678_ VGND net1320 net387 sg13g2_o21ai_1
XFILLER_33_990 VPWR VGND sg13g2_decap_8
X_4899_ _0615_ net1136 _0579_ _0616_ VPWR VGND sg13g2_a21o_1
X_3919_ _2299_ net928 _2298_ VPWR VGND sg13g2_nand2_1
XFILLER_3_349 VPWR VGND sg13g2_decap_4
Xfanout1117 net1118 net1117 VPWR VGND sg13g2_buf_8
Xfanout1128 net1129 net1128 VPWR VGND sg13g2_buf_8
Xfanout1106 net1107 net1106 VPWR VGND sg13g2_buf_2
XFILLER_47_504 VPWR VGND sg13g2_decap_8
XFILLER_47_21 VPWR VGND sg13g2_decap_8
Xfanout1139 net1140 net1139 VPWR VGND sg13g2_buf_8
XFILLER_15_401 VPWR VGND sg13g2_fill_2
XFILLER_28_795 VPWR VGND sg13g2_decap_8
XFILLER_16_968 VPWR VGND sg13g2_fill_2
XFILLER_16_979 VPWR VGND sg13g2_decap_8
XFILLER_7_600 VPWR VGND sg13g2_fill_1
XFILLER_6_110 VPWR VGND sg13g2_decap_4
XFILLER_12_90 VPWR VGND sg13g2_fill_1
XFILLER_40_7 VPWR VGND sg13g2_fill_1
XFILLER_3_894 VPWR VGND sg13g2_decap_8
X_5940_ _1553_ net1017 _1528_ _1554_ VPWR VGND sg13g2_a21o_1
XFILLER_19_795 VPWR VGND sg13g2_fill_2
X_5871_ _1491_ net467 net1031 VPWR VGND sg13g2_nand2b_1
X_4822_ net1149 VPWR _0546_ VGND _0544_ _0545_ sg13g2_o21ai_1
XFILLER_33_275 VPWR VGND sg13g2_fill_1
X_4753_ _0481_ net1144 _0430_ _0482_ VPWR VGND sg13g2_a21o_1
X_3704_ _2103_ net491 net977 VPWR VGND sg13g2_nand2b_1
X_4684_ s0.data_out\[16\]\[0\] s0.data_out\[17\]\[0\] net1164 _0421_ VPWR VGND sg13g2_mux2_1
X_3635_ _2037_ _2042_ _2043_ _2044_ VPWR VGND sg13g2_nor3_1
XFILLER_1_809 VPWR VGND sg13g2_decap_8
X_3566_ VPWR _0218_ net444 VGND sg13g2_inv_1
X_3497_ VGND VPWR _1856_ _1917_ _1918_ net1258 sg13g2_a21oi_1
XFILLER_0_308 VPWR VGND sg13g2_decap_8
X_5305_ VGND VPWR net1117 _0985_ _0986_ _0924_ sg13g2_a21oi_1
X_5236_ _0917_ _0920_ net1334 _0921_ VPWR VGND sg13g2_nand3_1
X_5167_ VGND VPWR net1129 _0859_ _0860_ _0800_ sg13g2_a21oi_1
X_5098_ net1127 VPWR _0796_ VGND _0794_ _0795_ sg13g2_o21ai_1
X_4118_ VPWR _2477_ net359 VGND sg13g2_inv_1
XFILLER_44_529 VPWR VGND sg13g2_decap_8
XFILLER_25_710 VPWR VGND sg13g2_fill_2
X_4049_ _2413_ VPWR _2414_ VGND _2465_ net1057 sg13g2_o21ai_1
XFILLER_17_68 VPWR VGND sg13g2_decap_8
XFILLER_13_949 VPWR VGND sg13g2_decap_8
XFILLER_3_124 VPWR VGND sg13g2_decap_4
XFILLER_3_168 VPWR VGND sg13g2_decap_8
XFILLER_0_831 VPWR VGND sg13g2_decap_8
Xhold8 s0.genblk1\[18\].modules.bubble VPWR VGND net304 sg13g2_dlygate4sd3_1
XFILLER_48_857 VPWR VGND sg13g2_decap_8
XFILLER_47_334 VPWR VGND sg13g2_fill_1
XFILLER_35_507 VPWR VGND sg13g2_decap_8
XFILLER_15_253 VPWR VGND sg13g2_decap_8
X_6207__273 VPWR VGND net273 sg13g2_tiehi
XFILLER_31_746 VPWR VGND sg13g2_fill_2
XFILLER_12_971 VPWR VGND sg13g2_decap_8
XFILLER_30_267 VPWR VGND sg13g2_fill_1
XFILLER_8_964 VPWR VGND sg13g2_decap_8
XFILLER_7_430 VPWR VGND sg13g2_decap_4
XFILLER_48_1011 VPWR VGND sg13g2_decap_8
X_3420_ _1846_ VPWR _1847_ VGND _1842_ _1845_ sg13g2_o21ai_1
X_3351_ _1734_ _1783_ _1784_ VPWR VGND sg13g2_and2_1
X_6070_ net210 VGND VPWR _0120_ s0.genblk1\[11\].modules.bubble clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
X_3282_ VGND VPWR net991 net463 _1722_ _1721_ sg13g2_a21oi_1
X_5021_ _0673_ _0725_ _0726_ VPWR VGND sg13g2_and2_1
XFILLER_38_334 VPWR VGND sg13g2_fill_2
XFILLER_0_1013 VPWR VGND sg13g2_decap_8
X_5923_ s0.data_out\[8\]\[1\] s0.data_out\[7\]\[1\] net1022 _1537_ VPWR VGND sg13g2_mux2_1
X_5854_ net1221 _1471_ _0165_ VPWR VGND sg13g2_nor2_1
XFILLER_34_584 VPWR VGND sg13g2_decap_8
X_4805_ net923 VPWR _0532_ VGND s0.was_valid_out\[15\][0] net1153 sg13g2_o21ai_1
XFILLER_22_746 VPWR VGND sg13g2_fill_1
XFILLER_22_757 VPWR VGND sg13g2_fill_2
XFILLER_22_768 VPWR VGND sg13g2_fill_1
X_5785_ VGND VPWR _1412_ net565 net1346 sg13g2_or2_1
X_4736_ net1305 VPWR _0467_ VGND _2462_ _0466_ sg13g2_o21ai_1
X_4667_ _0392_ _0407_ _0408_ VPWR VGND sg13g2_nor2b_1
X_3618_ VGND VPWR net983 _2026_ _2027_ _1987_ sg13g2_a21oi_1
XFILLER_1_606 VPWR VGND sg13g2_decap_8
X_4598_ VGND VPWR net1159 s0.data_out\[17\]\[5\] _0342_ _0341_ sg13g2_a21oi_1
X_6039__243 VPWR VGND net243 sg13g2_tiehi
X_3549_ _1963_ VPWR _1964_ VGND _1959_ _1962_ sg13g2_o21ai_1
X_6199_ net70 VGND VPWR _0249_ s0.valid_out\[1\][0] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_5219_ net1117 VPWR _0906_ VGND _0904_ _0905_ sg13g2_o21ai_1
XFILLER_28_45 VPWR VGND sg13g2_decap_4
XFILLER_29_334 VPWR VGND sg13g2_fill_1
XFILLER_29_345 VPWR VGND sg13g2_fill_2
XFILLER_45_816 VPWR VGND sg13g2_decap_8
XFILLER_44_348 VPWR VGND sg13g2_decap_8
X_6046__236 VPWR VGND net236 sg13g2_tiehi
XFILLER_25_562 VPWR VGND sg13g2_decap_8
XFILLER_8_205 VPWR VGND sg13g2_fill_2
XFILLER_5_923 VPWR VGND sg13g2_decap_8
XFILLER_48_654 VPWR VGND sg13g2_decap_8
XFILLER_47_120 VPWR VGND sg13g2_fill_2
XFILLER_47_164 VPWR VGND sg13g2_fill_1
XFILLER_47_153 VPWR VGND sg13g2_fill_1
XFILLER_44_871 VPWR VGND sg13g2_decap_8
XFILLER_12_790 VPWR VGND sg13g2_fill_2
X_5570_ _1119_ _1225_ _1226_ _1227_ VPWR VGND sg13g2_nor3_1
X_4521_ _0274_ net1176 net570 VPWR VGND sg13g2_nand2_1
Xhold216 _1992_ VPWR VGND net512 sg13g2_dlygate4sd3_1
X_4452_ net1287 VPWR _2773_ VGND net926 _2772_ sg13g2_o21ai_1
Xhold205 s0.data_out\[12\]\[5\] VPWR VGND net501 sg13g2_dlygate4sd3_1
Xhold249 _1642_ VPWR VGND net545 sg13g2_dlygate4sd3_1
Xhold227 s0.data_out\[20\]\[7\] VPWR VGND net523 sg13g2_dlygate4sd3_1
X_3403_ _1828_ _1831_ net1311 _1832_ VPWR VGND sg13g2_nand3_1
Xhold238 _1964_ VPWR VGND net534 sg13g2_dlygate4sd3_1
X_4383_ _2710_ net1180 _2684_ _2711_ VPWR VGND sg13g2_a21o_1
X_6122_ net154 VGND VPWR _0172_ s0.data_out\[8\]\[6\] clknet_leaf_17_clk sg13g2_dfrbpq_2
X_3334_ VPWR _0197_ net520 VGND sg13g2_inv_1
X_3265_ _2469_ VPWR _1708_ VGND net383 net1009 sg13g2_o21ai_1
X_6053_ net228 VGND VPWR _0103_ s0.data_out\[13\]\[4\] clknet_leaf_25_clk sg13g2_dfrbpq_2
X_5004_ VGND VPWR net1123 _0708_ _0709_ _0668_ sg13g2_a21oi_1
X_3196_ VPWR _0184_ net545 VGND sg13g2_inv_1
XFILLER_26_337 VPWR VGND sg13g2_decap_8
X_5906_ VGND VPWR net1017 net544 _1522_ _1521_ sg13g2_a21oi_1
XFILLER_22_521 VPWR VGND sg13g2_decap_8
X_5837_ _1460_ _1461_ _1462_ _1463_ VPWR VGND sg13g2_nor3_1
X_5768_ net1037 VPWR _1397_ VGND _1395_ _1396_ sg13g2_o21ai_1
X_4719_ net1146 net1057 _0452_ VPWR VGND sg13g2_nor2b_1
X_5699_ VGND VPWR _1344_ net1210 net315 sg13g2_or2_1
XFILLER_2_959 VPWR VGND sg13g2_decap_8
XFILLER_1_436 VPWR VGND sg13g2_decap_8
XFILLER_49_429 VPWR VGND sg13g2_decap_8
XFILLER_38_1010 VPWR VGND sg13g2_decap_8
XFILLER_40_351 VPWR VGND sg13g2_fill_2
XFILLER_20_90 VPWR VGND sg13g2_decap_8
XFILLER_1_970 VPWR VGND sg13g2_decap_8
XFILLER_49_996 VPWR VGND sg13g2_decap_8
XFILLER_36_635 VPWR VGND sg13g2_fill_1
XFILLER_24_819 VPWR VGND sg13g2_fill_2
XFILLER_35_167 VPWR VGND sg13g2_fill_1
X_3952_ net944 s0.data_out\[0\]\[5\] _2328_ VPWR VGND sg13g2_and2_1
X_3883_ VGND VPWR _2268_ _2267_ net1214 sg13g2_or2_1
X_5622_ net1082 VPWR _1271_ VGND _1269_ _1270_ sg13g2_o21ai_1
XFILLER_32_896 VPWR VGND sg13g2_fill_1
X_5553_ _1208_ _1209_ _1207_ _1210_ VPWR VGND sg13g2_nand3_1
X_4504_ _2819_ net1167 _2771_ _2820_ VPWR VGND sg13g2_a21o_1
X_5484_ _1146_ net436 net1096 VPWR VGND sg13g2_nand2b_1
X_4435_ net1167 net1069 _2758_ VPWR VGND sg13g2_nor2b_1
X_6216__136 VPWR VGND net136 sg13g2_tiehi
X_4366_ s0.data_out\[20\]\[1\] s0.data_out\[19\]\[1\] net1186 _2694_ VPWR VGND sg13g2_mux2_1
X_3317_ _1752_ VPWR _1753_ VGND _1748_ _1751_ sg13g2_o21ai_1
X_6036__246 VPWR VGND net246 sg13g2_tiehi
X_6105_ net172 VGND VPWR _0155_ s0.data_out\[9\]\[1\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_4297_ s0.data_out\[19\]\[0\] s0.data_out\[20\]\[0\] net1199 _2633_ VPWR VGND sg13g2_mux2_1
X_3248_ net1235 _1686_ _1693_ VPWR VGND sg13g2_nor2_1
X_6036_ net246 VGND VPWR _0086_ s0.valid_out\[14\][0] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_3179_ _1627_ VPWR _1628_ VGND _1623_ _1626_ sg13g2_o21ai_1
XFILLER_26_178 VPWR VGND sg13g2_decap_8
XFILLER_26_189 VPWR VGND sg13g2_fill_1
X_6043__239 VPWR VGND net239 sg13g2_tiehi
XFILLER_6_528 VPWR VGND sg13g2_fill_1
XFILLER_29_1009 VPWR VGND sg13g2_decap_8
XFILLER_2_756 VPWR VGND sg13g2_decap_8
XFILLER_49_259 VPWR VGND sg13g2_decap_8
XFILLER_46_922 VPWR VGND sg13g2_decap_8
XFILLER_46_999 VPWR VGND sg13g2_decap_8
XFILLER_14_841 VPWR VGND sg13g2_decap_4
XFILLER_32_115 VPWR VGND sg13g2_fill_1
XFILLER_14_852 VPWR VGND sg13g2_fill_1
XFILLER_32_148 VPWR VGND sg13g2_fill_2
XFILLER_9_311 VPWR VGND sg13g2_fill_2
XFILLER_9_366 VPWR VGND sg13g2_fill_1
XFILLER_12_1013 VPWR VGND sg13g2_decap_8
X_4220_ net1216 _2561_ _2562_ VPWR VGND sg13g2_nor2_1
X_4151_ _2502_ VPWR net9 VGND _2472_ net912 sg13g2_o21ai_1
X_4082_ net1342 net314 _0271_ VPWR VGND sg13g2_and2_1
XFILLER_49_793 VPWR VGND sg13g2_decap_8
XFILLER_37_999 VPWR VGND sg13g2_decap_8
XFILLER_24_605 VPWR VGND sg13g2_decap_4
X_4984_ _0691_ VPWR _0692_ VGND net1319 net438 sg13g2_o21ai_1
XFILLER_23_159 VPWR VGND sg13g2_decap_8
X_3935_ VGND VPWR _2245_ _2312_ _2313_ net951 sg13g2_a21oi_1
XFILLER_20_833 VPWR VGND sg13g2_fill_2
XFILLER_32_682 VPWR VGND sg13g2_fill_1
X_3866_ _2250_ VPWR _2251_ VGND _2243_ _2244_ sg13g2_o21ai_1
X_5605_ VGND VPWR net1040 net451 _1256_ _1255_ sg13g2_a21oi_1
X_3797_ _2188_ VPWR _2189_ VGND net1297 net426 sg13g2_o21ai_1
X_5536_ VPWR VGND _1126_ net1283 _1191_ net1278 _1193_ _1188_ sg13g2_a221oi_1
X_5467_ VPWR _0123_ _1131_ VGND sg13g2_inv_1
X_4418_ net1172 _2739_ _2744_ VPWR VGND sg13g2_nor2_1
X_5398_ _1067_ net1099 net536 VPWR VGND sg13g2_nand2_1
X_4349_ net1286 VPWR _2679_ VGND _2456_ _2678_ sg13g2_o21ai_1
XFILLER_46_218 VPWR VGND sg13g2_fill_2
X_6019_ net265 VGND VPWR _0069_ s0.data_out\[16\]\[6\] clknet_leaf_33_clk sg13g2_dfrbpq_2
XFILLER_27_454 VPWR VGND sg13g2_decap_8
XFILLER_43_947 VPWR VGND sg13g2_decap_8
XFILLER_14_137 VPWR VGND sg13g2_fill_2
XFILLER_35_1013 VPWR VGND sg13g2_decap_8
XFILLER_14_148 VPWR VGND sg13g2_fill_2
XFILLER_11_833 VPWR VGND sg13g2_fill_1
XFILLER_10_332 VPWR VGND sg13g2_fill_2
XFILLER_11_866 VPWR VGND sg13g2_fill_2
XFILLER_6_325 VPWR VGND sg13g2_decap_4
XFILLER_10_398 VPWR VGND sg13g2_fill_1
XFILLER_2_542 VPWR VGND sg13g2_decap_8
XFILLER_42_1006 VPWR VGND sg13g2_decap_8
XFILLER_2_586 VPWR VGND sg13g2_decap_4
XFILLER_37_207 VPWR VGND sg13g2_decap_8
XFILLER_19_966 VPWR VGND sg13g2_decap_8
XFILLER_46_796 VPWR VGND sg13g2_decap_8
XFILLER_18_487 VPWR VGND sg13g2_fill_2
XFILLER_33_402 VPWR VGND sg13g2_fill_1
X_3720_ _2117_ net968 net488 VPWR VGND sg13g2_nand2_1
X_3651_ net933 VPWR _2058_ VGND s0.was_valid_out\[2\][0] net977 sg13g2_o21ai_1
X_3582_ VPWR _0220_ net512 VGND sg13g2_inv_1
X_5321_ _0999_ VPWR _1000_ VGND net1105 _0879_ sg13g2_o21ai_1
X_5252_ VGND VPWR _0935_ net597 net1338 sg13g2_or2_1
X_5183_ _0765_ _0874_ _0875_ _0876_ VPWR VGND sg13g2_nor3_1
X_4203_ net1205 _2545_ _2546_ _2547_ VPWR VGND sg13g2_nor3_1
XFILLER_29_719 VPWR VGND sg13g2_decap_8
X_4134_ VPWR _2493_ s0.data_out\[1\]\[2\] VGND sg13g2_inv_1
XFILLER_49_590 VPWR VGND sg13g2_decap_8
X_4065_ VGND VPWR _2426_ _2419_ net1246 sg13g2_or2_1
XFILLER_25_914 VPWR VGND sg13g2_fill_2
XFILLER_19_1008 VPWR VGND sg13g2_decap_8
XFILLER_24_468 VPWR VGND sg13g2_decap_8
XFILLER_24_479 VPWR VGND sg13g2_fill_2
X_4967_ _0677_ _0673_ _0676_ VPWR VGND sg13g2_nand2b_1
Xclkbuf_leaf_31_clk clknet_3_4__leaf_clk clknet_leaf_31_clk VPWR VGND sg13g2_buf_8
X_4898_ s0.data_out\[16\]\[6\] s0.data_out\[15\]\[6\] net1143 _0615_ VPWR VGND sg13g2_mux2_1
X_3918_ s0.data_out\[0\]\[1\] s0.data_out\[1\]\[1\] net955 _2298_ VPWR VGND sg13g2_mux2_1
XFILLER_32_490 VPWR VGND sg13g2_decap_8
XFILLER_22_58 VPWR VGND sg13g2_decap_8
X_3849_ VGND VPWR net961 _2233_ _2234_ _2191_ sg13g2_a21oi_1
X_5519_ VGND VPWR net1080 net531 _1177_ _1176_ sg13g2_a21oi_1
XFILLER_0_7 VPWR VGND sg13g2_decap_8
Xfanout1118 s0.shift_out\[13\][0] net1118 VPWR VGND sg13g2_buf_8
Xfanout1129 net335 net1129 VPWR VGND sg13g2_buf_8
Xfanout1107 s0.shift_out\[12\][0] net1107 VPWR VGND sg13g2_buf_8
XFILLER_47_527 VPWR VGND sg13g2_decap_8
XFILLER_42_254 VPWR VGND sg13g2_fill_2
XFILLER_42_232 VPWR VGND sg13g2_fill_2
XFILLER_15_446 VPWR VGND sg13g2_decap_4
XFILLER_8_49 VPWR VGND sg13g2_decap_4
XFILLER_8_16 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_22_clk clknet_3_6__leaf_clk clknet_leaf_22_clk VPWR VGND sg13g2_buf_8
XFILLER_7_634 VPWR VGND sg13g2_fill_1
XFILLER_10_173 VPWR VGND sg13g2_decap_4
XFILLER_3_873 VPWR VGND sg13g2_decap_8
XFILLER_2_350 VPWR VGND sg13g2_fill_1
XFILLER_2_394 VPWR VGND sg13g2_fill_2
X_5870_ VPWR _0167_ _1490_ VGND sg13g2_inv_1
X_4821_ net1135 net1070 _0545_ VPWR VGND sg13g2_nor2b_1
XFILLER_15_980 VPWR VGND sg13g2_decap_8
XFILLER_21_405 VPWR VGND sg13g2_decap_8
XFILLER_33_287 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_13_clk clknet_3_3__leaf_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
X_4752_ s0.data_out\[17\]\[1\] s0.data_out\[16\]\[1\] net1151 _0481_ VPWR VGND sg13g2_mux2_1
XFILLER_33_298 VPWR VGND sg13g2_decap_4
X_3703_ VPWR _0231_ _2102_ VGND sg13g2_inv_1
X_4683_ net1219 _0419_ _0050_ VPWR VGND sg13g2_nor2_1
X_3634_ VGND VPWR _1980_ _2035_ _2043_ net1249 sg13g2_a21oi_1
X_3565_ _1977_ VPWR _1978_ VGND net1308 net443 sg13g2_o21ai_1
X_3496_ _1917_ net993 _1916_ VPWR VGND sg13g2_nand2b_1
X_5304_ _0984_ net1106 _0925_ _0985_ VPWR VGND sg13g2_a21o_1
X_5235_ net1116 VPWR _0920_ VGND _0918_ _0919_ sg13g2_o21ai_1
X_5166_ _0858_ net1115 _0801_ _0859_ VPWR VGND sg13g2_a21o_1
X_5097_ net1113 net1063 _0795_ VPWR VGND sg13g2_nor2b_1
X_4117_ VPWR _2476_ net1254 VGND sg13g2_inv_1
XFILLER_44_519 VPWR VGND sg13g2_fill_1
X_4048_ net374 net946 net941 _2413_ VPWR VGND sg13g2_a21o_1
XFILLER_25_733 VPWR VGND sg13g2_decap_8
XFILLER_13_917 VPWR VGND sg13g2_decap_8
XFILLER_24_221 VPWR VGND sg13g2_fill_1
XFILLER_13_928 VPWR VGND sg13g2_decap_8
X_5999_ net287 VGND VPWR net376 s0.was_valid_out\[17\][0] clknet_leaf_33_clk sg13g2_dfrbpq_1
XFILLER_21_983 VPWR VGND sg13g2_decap_8
XFILLER_20_471 VPWR VGND sg13g2_fill_2
XFILLER_4_637 VPWR VGND sg13g2_fill_2
XFILLER_0_810 VPWR VGND sg13g2_decap_8
X_5994__292 VPWR VGND net292 sg13g2_tiehi
XFILLER_48_836 VPWR VGND sg13g2_decap_8
XFILLER_0_887 VPWR VGND sg13g2_decap_8
Xhold9 s0.genblk1\[19\].modules.bubble VPWR VGND net305 sg13g2_dlygate4sd3_1
XFILLER_47_379 VPWR VGND sg13g2_fill_1
XFILLER_16_722 VPWR VGND sg13g2_decap_8
XFILLER_16_733 VPWR VGND sg13g2_decap_4
XFILLER_15_232 VPWR VGND sg13g2_decap_8
XFILLER_12_950 VPWR VGND sg13g2_decap_8
XFILLER_8_943 VPWR VGND sg13g2_decap_8
X_3350_ _1783_ net1003 _1782_ VPWR VGND sg13g2_nand2b_1
X_5020_ _0725_ net1138 _0724_ VPWR VGND sg13g2_nand2b_1
X_3281_ net992 net1070 _1721_ VPWR VGND sg13g2_nor2b_1
XFILLER_31_4 VPWR VGND sg13g2_fill_1
XFILLER_39_814 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_2_clk clknet_3_0__leaf_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
XFILLER_17_2 VPWR VGND sg13g2_fill_1
XFILLER_26_508 VPWR VGND sg13g2_decap_8
XFILLER_26_519 VPWR VGND sg13g2_fill_2
XFILLER_19_582 VPWR VGND sg13g2_fill_1
XFILLER_0_83 VPWR VGND sg13g2_decap_8
X_5922_ VGND VPWR _1536_ _1535_ net1272 sg13g2_or2_1
X_5853_ VGND VPWR _1472_ _1475_ _0164_ _1476_ sg13g2_a21oi_1
XFILLER_21_202 VPWR VGND sg13g2_decap_8
XFILLER_22_714 VPWR VGND sg13g2_fill_1
X_5784_ net1343 VPWR _1411_ VGND net920 _1410_ sg13g2_o21ai_1
X_4804_ net1136 _0525_ _0531_ VPWR VGND sg13g2_nor2_1
XFILLER_21_235 VPWR VGND sg13g2_fill_1
XFILLER_9_70 VPWR VGND sg13g2_decap_4
X_4735_ VGND VPWR net1146 net546 _0466_ _0465_ sg13g2_a21oi_1
X_4666_ _0397_ VPWR _0407_ VGND _0403_ _0404_ sg13g2_o21ai_1
X_3617_ _2025_ net972 _1988_ _2026_ VPWR VGND sg13g2_a21o_1
X_4597_ net1159 net1054 _0341_ VPWR VGND sg13g2_nor2b_1
X_3548_ VGND VPWR _1963_ net533 net1312 sg13g2_or2_1
X_3479_ _1849_ _1899_ _1900_ VPWR VGND sg13g2_and2_1
X_6198_ net72 VGND VPWR net329 s0.was_valid_out\[1\][0] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_5218_ net1101 net1066 _0905_ VPWR VGND sg13g2_nor2b_1
X_5149_ VGND VPWR net1113 _0841_ _0842_ _0795_ sg13g2_a21oi_1
XFILLER_40_511 VPWR VGND sg13g2_fill_1
XFILLER_40_544 VPWR VGND sg13g2_fill_2
XFILLER_40_566 VPWR VGND sg13g2_fill_1
XFILLER_5_902 VPWR VGND sg13g2_decap_8
XFILLER_4_401 VPWR VGND sg13g2_fill_2
XFILLER_5_979 VPWR VGND sg13g2_decap_8
XFILLER_4_467 VPWR VGND sg13g2_fill_1
XFILLER_48_633 VPWR VGND sg13g2_decap_8
XFILLER_0_684 VPWR VGND sg13g2_decap_8
XFILLER_10_9 VPWR VGND sg13g2_decap_4
XFILLER_44_850 VPWR VGND sg13g2_decap_8
XFILLER_16_585 VPWR VGND sg13g2_decap_8
XFILLER_15_1022 VPWR VGND sg13g2_decap_8
X_4520_ _0272_ _2833_ _0273_ VPWR VGND _2834_ sg13g2_nand3b_1
X_4451_ VGND VPWR net1167 net478 _2772_ _2771_ sg13g2_a21oi_1
Xhold206 _1047_ VPWR VGND net502 sg13g2_dlygate4sd3_1
Xhold217 s0.data_out\[1\]\[3\] VPWR VGND net513 sg13g2_dlygate4sd3_1
Xhold239 s0.data_out\[4\]\[7\] VPWR VGND net535 sg13g2_dlygate4sd3_1
Xhold228 _2688_ VPWR VGND net524 sg13g2_dlygate4sd3_1
X_3402_ net990 VPWR _1831_ VGND _1829_ _1830_ sg13g2_o21ai_1
X_6121_ net155 VGND VPWR _0171_ s0.data_out\[8\]\[5\] clknet_leaf_18_clk sg13g2_dfrbpq_2
X_4382_ s0.data_out\[20\]\[7\] s0.data_out\[19\]\[7\] net1186 _2710_ VPWR VGND sg13g2_mux2_1
X_3333_ _1766_ VPWR _1767_ VGND _1762_ _1765_ sg13g2_o21ai_1
X_3264_ VGND VPWR _1707_ net999 net383 sg13g2_or2_1
X_6052_ net229 VGND VPWR _0102_ s0.data_out\[13\]\[3\] clknet_leaf_29_clk sg13g2_dfrbpq_2
XFILLER_39_622 VPWR VGND sg13g2_fill_1
XFILLER_38_121 VPWR VGND sg13g2_fill_2
X_5003_ s0.data_out\[15\]\[2\] s0.data_out\[14\]\[2\] net1130 _0708_ VPWR VGND sg13g2_mux2_1
X_3195_ _1641_ VPWR _1642_ VGND _1637_ _1640_ sg13g2_o21ai_1
XFILLER_38_154 VPWR VGND sg13g2_fill_1
Xfanout1290 net1291 net1290 VPWR VGND sg13g2_buf_8
XFILLER_27_806 VPWR VGND sg13g2_decap_8
XFILLER_27_817 VPWR VGND sg13g2_fill_1
X_5905_ net1017 net1051 _1521_ VPWR VGND sg13g2_nor2b_1
XFILLER_34_382 VPWR VGND sg13g2_fill_1
X_5836_ VGND VPWR _1387_ _1457_ _1462_ net1257 sg13g2_a21oi_1
XFILLER_22_577 VPWR VGND sg13g2_fill_2
X_5767_ net1027 net1055 _1396_ VPWR VGND sg13g2_nor2b_1
X_4718_ net1146 s0.data_out\[16\]\[4\] _0451_ VPWR VGND sg13g2_and2_1
X_6178__93 VPWR VGND net93 sg13g2_tiehi
XFILLER_30_14 VPWR VGND sg13g2_decap_8
X_5698_ VPWR VGND _1342_ _1233_ _1327_ _1323_ _1343_ _1325_ sg13g2_a221oi_1
X_4649_ net1240 _0388_ _0390_ VPWR VGND sg13g2_nor2_1
XFILLER_2_938 VPWR VGND sg13g2_decap_8
XFILLER_49_408 VPWR VGND sg13g2_decap_8
XFILLER_45_614 VPWR VGND sg13g2_fill_1
XFILLER_45_1026 VPWR VGND sg13g2_fill_2
XFILLER_49_975 VPWR VGND sg13g2_decap_8
XFILLER_48_485 VPWR VGND sg13g2_decap_8
X_3951_ _2327_ net929 _2326_ VPWR VGND sg13g2_nand2_1
XFILLER_16_393 VPWR VGND sg13g2_fill_2
X_3882_ _2205_ VPWR _2267_ VGND net930 _2266_ sg13g2_o21ai_1
X_6029__254 VPWR VGND net254 sg13g2_tiehi
X_5621_ net1040 net1060 _1270_ VPWR VGND sg13g2_nor2b_1
X_5552_ VGND VPWR _1209_ _1202_ net1237 sg13g2_or2_1
X_4503_ s0.data_out\[19\]\[3\] s0.data_out\[18\]\[3\] net1174 _2819_ VPWR VGND sg13g2_mux2_1
X_6175__96 VPWR VGND net96 sg13g2_tiehi
X_5483_ VPWR _0125_ _1145_ VGND sg13g2_inv_1
X_4434_ net925 _2484_ _2757_ VPWR VGND sg13g2_nor2_1
X_4365_ _2693_ net1187 s0.data_out\[19\]\[1\] VPWR VGND sg13g2_nand2_1
X_3316_ VGND VPWR _1752_ net539 net1325 sg13g2_or2_1
X_6104_ net173 VGND VPWR _0154_ s0.data_out\[9\]\[0\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_6035_ net248 VGND VPWR _0085_ s0.was_valid_out\[14\][0] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_4296_ net1217 _2626_ _0014_ VPWR VGND sg13g2_nor2_1
XFILLER_39_452 VPWR VGND sg13g2_decap_4
XFILLER_39_430 VPWR VGND sg13g2_fill_2
X_3247_ VGND VPWR _1692_ _1690_ net1244 sg13g2_or2_1
X_3178_ VGND VPWR _1627_ net411 net1329 sg13g2_or2_1
XFILLER_27_625 VPWR VGND sg13g2_fill_1
XFILLER_42_628 VPWR VGND sg13g2_fill_1
XFILLER_25_25 VPWR VGND sg13g2_decap_8
XFILLER_23_842 VPWR VGND sg13g2_decap_8
X_5819_ VPWR _1445_ _1444_ VGND sg13g2_inv_1
XFILLER_10_514 VPWR VGND sg13g2_decap_8
XFILLER_6_507 VPWR VGND sg13g2_decap_8
XFILLER_2_735 VPWR VGND sg13g2_decap_8
XFILLER_49_227 VPWR VGND sg13g2_decap_8
XFILLER_46_901 VPWR VGND sg13g2_decap_8
XFILLER_18_625 VPWR VGND sg13g2_decap_8
XFILLER_46_978 VPWR VGND sg13g2_decap_8
XFILLER_45_422 VPWR VGND sg13g2_fill_1
XFILLER_14_864 VPWR VGND sg13g2_fill_1
XFILLER_40_171 VPWR VGND sg13g2_fill_1
XFILLER_9_334 VPWR VGND sg13g2_fill_1
XFILLER_40_193 VPWR VGND sg13g2_decap_8
XFILLER_40_182 VPWR VGND sg13g2_fill_1
XFILLER_9_389 VPWR VGND sg13g2_decap_8
X_4150_ _2502_ net1231 _2494_ VPWR VGND sg13g2_nand2_1
X_4081_ _2440_ _2441_ _0270_ VPWR VGND sg13g2_and2_1
XFILLER_49_772 VPWR VGND sg13g2_decap_8
XFILLER_37_978 VPWR VGND sg13g2_decap_8
XFILLER_36_422 VPWR VGND sg13g2_fill_2
XFILLER_24_617 VPWR VGND sg13g2_decap_8
XFILLER_17_680 VPWR VGND sg13g2_fill_1
X_4983_ _0687_ _0690_ net1323 _0691_ VPWR VGND sg13g2_nand3_1
X_3934_ _2312_ net348 net955 VPWR VGND sg13g2_nand2b_1
X_3865_ _2250_ _2249_ net1261 _2234_ net1268 VPWR VGND sg13g2_a22oi_1
X_5604_ net1040 net1067 _1255_ VPWR VGND sg13g2_nor2b_1
X_6042__240 VPWR VGND net240 sg13g2_tiehi
XFILLER_20_889 VPWR VGND sg13g2_fill_1
X_3796_ _2184_ _2187_ net1297 _2188_ VPWR VGND sg13g2_nand3_1
X_5535_ net1278 _1188_ _1192_ VPWR VGND sg13g2_nor2_1
X_5466_ _1130_ VPWR _1131_ VGND net1335 net452 sg13g2_o21ai_1
X_4417_ _2741_ VPWR _2743_ VGND s0.was_valid_out\[18\][0] net1176 sg13g2_o21ai_1
X_5397_ net1270 _1065_ _1066_ VPWR VGND sg13g2_nor2_1
XFILLER_28_1021 VPWR VGND sg13g2_decap_8
X_4348_ VGND VPWR net1182 net551 _2678_ _2677_ sg13g2_a21oi_1
X_4279_ _2602_ _2618_ _2619_ VPWR VGND sg13g2_nor2b_1
XFILLER_39_271 VPWR VGND sg13g2_fill_1
XFILLER_39_260 VPWR VGND sg13g2_decap_4
X_6018_ net266 VGND VPWR _0068_ s0.data_out\[16\]\[5\] clknet_leaf_32_clk sg13g2_dfrbpq_2
XFILLER_28_923 VPWR VGND sg13g2_decap_4
XFILLER_36_24 VPWR VGND sg13g2_decap_4
XFILLER_27_433 VPWR VGND sg13g2_decap_8
XFILLER_43_926 VPWR VGND sg13g2_decap_8
XFILLER_36_68 VPWR VGND sg13g2_fill_2
XFILLER_36_57 VPWR VGND sg13g2_decap_8
XFILLER_15_617 VPWR VGND sg13g2_fill_1
XFILLER_42_414 VPWR VGND sg13g2_fill_1
XFILLER_14_116 VPWR VGND sg13g2_decap_4
XFILLER_42_458 VPWR VGND sg13g2_fill_1
XFILLER_30_609 VPWR VGND sg13g2_decap_8
XFILLER_22_160 VPWR VGND sg13g2_decap_8
XFILLER_10_322 VPWR VGND sg13g2_fill_1
XFILLER_10_355 VPWR VGND sg13g2_fill_1
XFILLER_10_377 VPWR VGND sg13g2_decap_8
XFILLER_6_348 VPWR VGND sg13g2_decap_8
XFILLER_2_510 VPWR VGND sg13g2_fill_1
XFILLER_38_709 VPWR VGND sg13g2_fill_1
XFILLER_18_411 VPWR VGND sg13g2_fill_1
XFILLER_46_775 VPWR VGND sg13g2_decap_8
XFILLER_33_414 VPWR VGND sg13g2_decap_8
XFILLER_42_992 VPWR VGND sg13g2_decap_8
X_6026__257 VPWR VGND net257 sg13g2_tiehi
X_3650_ net963 _2051_ _2057_ VPWR VGND sg13g2_nor2_1
X_3581_ _1991_ VPWR _1992_ VGND _1987_ _1990_ sg13g2_o21ai_1
XFILLER_6_871 VPWR VGND sg13g2_fill_1
X_5320_ VPWR _0999_ _0998_ VGND sg13g2_inv_1
X_5251_ net1338 VPWR _0934_ VGND net936 _0933_ sg13g2_o21ai_1
X_4202_ net1207 s0.data_out\[20\]\[4\] _2546_ VPWR VGND sg13g2_nor2_1
X_5182_ _0854_ _0855_ _0875_ VPWR VGND sg13g2_nor2b_1
X_4133_ VPWR _2492_ s0.data_out\[3\]\[2\] VGND sg13g2_inv_1
X_4064_ VGND VPWR net1294 _2425_ _0269_ _2423_ sg13g2_a21oi_1
XFILLER_25_926 VPWR VGND sg13g2_decap_4
X_4966_ net1320 VPWR _0676_ VGND net921 _0675_ sg13g2_o21ai_1
X_4897_ _0614_ net1142 net562 VPWR VGND sg13g2_nand2_1
X_3917_ VPWR _0250_ net449 VGND sg13g2_inv_1
X_3848_ _2232_ net949 _2192_ _2233_ VPWR VGND sg13g2_a21o_1
X_3779_ VPWR _2174_ _2173_ VGND sg13g2_inv_1
XFILLER_20_697 VPWR VGND sg13g2_fill_1
X_5518_ net1080 net1047 _1176_ VPWR VGND sg13g2_nor2b_1
X_5449_ net1229 net1085 _1116_ VPWR VGND sg13g2_nor2b_1
Xfanout1119 net1120 net1119 VPWR VGND sg13g2_buf_8
Xfanout1108 s0.valid_out\[12\][0] net1108 VPWR VGND sg13g2_buf_8
XFILLER_19_208 VPWR VGND sg13g2_decap_4
XFILLER_19_219 VPWR VGND sg13g2_fill_1
XFILLER_28_720 VPWR VGND sg13g2_fill_1
XFILLER_42_200 VPWR VGND sg13g2_fill_1
XFILLER_42_222 VPWR VGND sg13g2_decap_4
XFILLER_23_480 VPWR VGND sg13g2_decap_8
XFILLER_11_675 VPWR VGND sg13g2_fill_2
XFILLER_7_679 VPWR VGND sg13g2_decap_8
XFILLER_12_81 VPWR VGND sg13g2_decap_8
XFILLER_3_852 VPWR VGND sg13g2_decap_8
XFILLER_19_753 VPWR VGND sg13g2_decap_8
X_6212__195 VPWR VGND net195 sg13g2_tiehi
XFILLER_19_797 VPWR VGND sg13g2_fill_1
X_4820_ net1135 s0.data_out\[15\]\[1\] _0544_ VPWR VGND sg13g2_and2_1
XFILLER_22_907 VPWR VGND sg13g2_decap_8
X_4751_ VGND VPWR _0480_ _0479_ net1268 sg13g2_or2_1
XFILLER_30_951 VPWR VGND sg13g2_fill_2
X_3702_ _2101_ VPWR _2102_ VGND _2097_ _2100_ sg13g2_o21ai_1
X_4682_ VGND VPWR _0415_ _0418_ _0049_ _0420_ sg13g2_a21oi_1
X_6220__84 VPWR VGND net84 sg13g2_tiehi
X_3633_ _2042_ net1215 _2040_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_995 VPWR VGND sg13g2_decap_8
X_3564_ _1973_ _1976_ net1308 _1977_ VPWR VGND sg13g2_nand3_1
X_3495_ VGND VPWR net982 _1915_ _1916_ _1858_ sg13g2_a21oi_1
X_5303_ s0.data_out\[13\]\[5\] s0.data_out\[12\]\[5\] net1110 _0984_ VPWR VGND sg13g2_mux2_1
X_5234_ net1102 net1060 _0919_ VPWR VGND sg13g2_nor2b_1
X_5165_ s0.data_out\[14\]\[4\] s0.data_out\[13\]\[4\] net1120 _0858_ VPWR VGND sg13g2_mux2_1
XFILLER_25_1013 VPWR VGND sg13g2_decap_8
X_4116_ VPWR _2475_ net361 VGND sg13g2_inv_1
XFILLER_29_506 VPWR VGND sg13g2_decap_4
X_5096_ net1113 s0.data_out\[13\]\[3\] _0794_ VPWR VGND sg13g2_and2_1
X_4047_ VGND VPWR net1292 _2412_ _0265_ _2410_ sg13g2_a21oi_1
XFILLER_37_572 VPWR VGND sg13g2_decap_4
XFILLER_25_712 VPWR VGND sg13g2_fill_1
XFILLER_40_737 VPWR VGND sg13g2_fill_2
X_5998_ net288 VGND VPWR _0048_ s0.genblk1\[17\].modules.bubble clknet_leaf_4_clk
+ sg13g2_dfrbpq_1
X_4949_ net1122 net1070 _0661_ VPWR VGND sg13g2_nor2b_1
XFILLER_24_288 VPWR VGND sg13g2_decap_8
XFILLER_32_1017 VPWR VGND sg13g2_decap_8
XFILLER_32_1028 VPWR VGND sg13g2_fill_1
XFILLER_20_483 VPWR VGND sg13g2_fill_2
XFILLER_4_649 VPWR VGND sg13g2_fill_1
XFILLER_0_866 VPWR VGND sg13g2_decap_8
XFILLER_48_815 VPWR VGND sg13g2_decap_8
XFILLER_47_347 VPWR VGND sg13g2_fill_2
XFILLER_15_211 VPWR VGND sg13g2_decap_4
XFILLER_30_203 VPWR VGND sg13g2_decap_4
XFILLER_8_922 VPWR VGND sg13g2_decap_8
XFILLER_8_900 VPWR VGND sg13g2_decap_4
XFILLER_7_476 VPWR VGND sg13g2_fill_1
XFILLER_7_454 VPWR VGND sg13g2_fill_2
XFILLER_8_999 VPWR VGND sg13g2_decap_8
X_3280_ VGND VPWR _1654_ _1719_ _1720_ net1000 sg13g2_a21oi_1
XFILLER_24_4 VPWR VGND sg13g2_fill_2
XFILLER_47_892 VPWR VGND sg13g2_decap_8
XFILLER_0_51 VPWR VGND sg13g2_fill_1
XFILLER_0_40 VPWR VGND sg13g2_decap_8
X_5921_ VGND VPWR net1023 _1534_ _1535_ _1492_ sg13g2_a21oi_1
X_5852_ net1342 VPWR _1476_ VGND net398 _1471_ sg13g2_o21ai_1
XFILLER_34_575 VPWR VGND sg13g2_decap_4
X_5783_ VGND VPWR net1028 s0.data_out\[8\]\[7\] _1410_ _1409_ sg13g2_a21oi_1
X_4803_ _0527_ VPWR _0530_ VGND s0.was_valid_out\[15\][0] net1141 sg13g2_o21ai_1
X_4734_ net1147 net1049 _0465_ VPWR VGND sg13g2_nor2b_1
X_4665_ _0402_ _0403_ _0380_ _0406_ VPWR VGND _0405_ sg13g2_nand4_1
X_3616_ s0.data_out\[4\]\[6\] s0.data_out\[3\]\[6\] net978 _2025_ VPWR VGND sg13g2_mux2_1
X_4596_ VGND VPWR _0274_ _0339_ _0340_ net1172 sg13g2_a21oi_1
X_3547_ net1312 VPWR _1962_ VGND net914 _1961_ sg13g2_o21ai_1
XFILLER_0_129 VPWR VGND sg13g2_decap_8
X_3478_ _1899_ net990 _1898_ VPWR VGND sg13g2_nand2b_1
X_5217_ net1100 net612 _0904_ VPWR VGND sg13g2_and2_1
X_6197_ net73 VGND VPWR _0247_ s0.genblk1\[21\].modules.bubble clknet_leaf_1_clk sg13g2_dfrbpq_1
X_5148_ _0840_ VPWR _0841_ VGND net1119 _2486_ sg13g2_o21ai_1
XFILLER_29_314 VPWR VGND sg13g2_decap_4
X_5079_ VGND VPWR _0712_ _0778_ _0779_ net1127 sg13g2_a21oi_1
XFILLER_44_35 VPWR VGND sg13g2_fill_1
XFILLER_13_726 VPWR VGND sg13g2_decap_8
XFILLER_40_578 VPWR VGND sg13g2_decap_8
XFILLER_8_207 VPWR VGND sg13g2_fill_1
XFILLER_20_280 VPWR VGND sg13g2_fill_1
XFILLER_5_958 VPWR VGND sg13g2_decap_8
XFILLER_4_413 VPWR VGND sg13g2_fill_2
XFILLER_48_612 VPWR VGND sg13g2_decap_8
XFILLER_0_663 VPWR VGND sg13g2_decap_8
XFILLER_47_111 VPWR VGND sg13g2_fill_1
XFILLER_48_689 VPWR VGND sg13g2_decap_8
XFILLER_29_881 VPWR VGND sg13g2_decap_8
XFILLER_35_339 VPWR VGND sg13g2_fill_1
XFILLER_43_383 VPWR VGND sg13g2_fill_2
XFILLER_15_1001 VPWR VGND sg13g2_decap_8
X_6187__83 VPWR VGND net83 sg13g2_tiehi
XFILLER_31_589 VPWR VGND sg13g2_decap_8
X_4450_ net1167 net1061 _2771_ VPWR VGND sg13g2_nor2b_1
Xhold207 s0.data_out\[7\]\[3\] VPWR VGND net503 sg13g2_dlygate4sd3_1
X_4381_ _2709_ net1186 net574 VPWR VGND sg13g2_nand2_1
Xhold229 s0.data_out\[14\]\[4\] VPWR VGND net525 sg13g2_dlygate4sd3_1
X_3401_ net981 net1074 _1830_ VPWR VGND sg13g2_nor2b_1
Xhold218 _2318_ VPWR VGND net514 sg13g2_dlygate4sd3_1
X_3332_ VGND VPWR _1766_ net519 net1325 sg13g2_or2_1
X_6120_ net156 VGND VPWR _0170_ s0.data_out\[8\]\[4\] clknet_leaf_18_clk sg13g2_dfrbpq_2
XFILLER_4_991 VPWR VGND sg13g2_decap_8
X_3263_ _1705_ VPWR _1706_ VGND net1004 _1585_ sg13g2_o21ai_1
X_6051_ net230 VGND VPWR _0101_ s0.data_out\[13\]\[2\] clknet_leaf_29_clk sg13g2_dfrbpq_2
X_3194_ VGND VPWR _1641_ net544 net1329 sg13g2_or2_1
X_5002_ _0707_ net1131 net573 VPWR VGND sg13g2_nand2_1
XFILLER_15_0 VPWR VGND sg13g2_fill_1
Xfanout1291 net1350 net1291 VPWR VGND sg13g2_buf_8
XFILLER_22_1027 VPWR VGND sg13g2_fill_2
Xfanout1280 ui_in[1] net1280 VPWR VGND sg13g2_buf_8
XFILLER_38_166 VPWR VGND sg13g2_fill_2
X_5904_ VGND VPWR _1440_ _1519_ _1520_ net1025 sg13g2_a21oi_1
XFILLER_35_873 VPWR VGND sg13g2_fill_1
Xclkbuf_3_5__f_clk clknet_0_clk clknet_3_5__leaf_clk VPWR VGND sg13g2_buf_8
X_5835_ net1266 _1432_ _1461_ VPWR VGND sg13g2_nor2_1
XFILLER_10_718 VPWR VGND sg13g2_decap_8
XFILLER_22_545 VPWR VGND sg13g2_fill_1
X_5766_ net1029 net610 _1395_ VPWR VGND sg13g2_and2_1
X_4717_ _0450_ net924 _0449_ VPWR VGND sg13g2_nand2_1
X_5697_ _1335_ VPWR _1342_ VGND _1331_ _1339_ sg13g2_o21ai_1
X_4648_ _0389_ _0388_ net1240 _0384_ net1233 VPWR VGND sg13g2_a22oi_1
X_4579_ s0.data_out\[17\]\[3\] s0.data_out\[18\]\[3\] net1175 _0325_ VPWR VGND sg13g2_mux2_1
XFILLER_2_917 VPWR VGND sg13g2_decap_8
XFILLER_29_133 VPWR VGND sg13g2_decap_8
XFILLER_29_188 VPWR VGND sg13g2_decap_8
XFILLER_44_125 VPWR VGND sg13g2_fill_2
XFILLER_41_843 VPWR VGND sg13g2_decap_4
XFILLER_41_876 VPWR VGND sg13g2_decap_8
XFILLER_40_353 VPWR VGND sg13g2_fill_1
XFILLER_9_516 VPWR VGND sg13g2_decap_8
XFILLER_41_898 VPWR VGND sg13g2_decap_8
XFILLER_20_70 VPWR VGND sg13g2_fill_2
XFILLER_45_1005 VPWR VGND sg13g2_decap_8
XFILLER_49_954 VPWR VGND sg13g2_decap_8
XFILLER_48_464 VPWR VGND sg13g2_decap_8
Xhold90 s0.data_out\[14\]\[3\] VPWR VGND net386 sg13g2_dlygate4sd3_1
X_6168__104 VPWR VGND net104 sg13g2_tiehi
XFILLER_35_103 VPWR VGND sg13g2_fill_2
X_3950_ s0.data_out\[0\]\[5\] s0.data_out\[1\]\[5\] net956 _2326_ VPWR VGND sg13g2_mux2_1
XFILLER_17_862 VPWR VGND sg13g2_decap_8
XFILLER_32_843 VPWR VGND sg13g2_decap_4
X_3881_ VGND VPWR net950 _2265_ _2266_ _2207_ sg13g2_a21oi_1
XFILLER_31_342 VPWR VGND sg13g2_fill_2
XFILLER_32_854 VPWR VGND sg13g2_decap_8
X_5620_ net1040 s0.data_out\[9\]\[4\] _1269_ VPWR VGND sg13g2_and2_1
X_5551_ VGND VPWR _1208_ _1206_ net1243 sg13g2_or2_1
X_4502_ VPWR VGND _2817_ _2813_ _2812_ net1212 _2818_ _2807_ sg13g2_a221oi_1
X_5482_ _1144_ VPWR _1145_ VGND _1140_ _1143_ sg13g2_o21ai_1
XFILLER_6_83 VPWR VGND sg13g2_decap_8
X_4433_ _2756_ net926 _2755_ VPWR VGND sg13g2_nand2_1
X_4364_ VGND VPWR _2692_ _2691_ net1268 sg13g2_or2_1
X_3315_ net1325 VPWR _1751_ VGND net916 _1750_ sg13g2_o21ai_1
X_6103_ net174 VGND VPWR _0153_ s0.valid_out\[9\][0] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_4295_ VGND VPWR _2628_ _2631_ _0013_ _2632_ sg13g2_a21oi_1
X_3246_ _1691_ _1690_ net1244 _1686_ net1235 VPWR VGND sg13g2_a22oi_1
XFILLER_6_1010 VPWR VGND sg13g2_decap_8
X_6034_ net249 VGND VPWR _0084_ s0.genblk1\[14\].modules.bubble clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
X_3177_ net1329 VPWR _1626_ VGND _2468_ _1625_ sg13g2_o21ai_1
XFILLER_35_670 VPWR VGND sg13g2_fill_2
XFILLER_23_865 VPWR VGND sg13g2_fill_2
X_5818_ _1444_ _1443_ net1243 _1439_ net1237 VPWR VGND sg13g2_a22oi_1
XFILLER_41_36 VPWR VGND sg13g2_fill_2
XFILLER_10_548 VPWR VGND sg13g2_fill_1
X_5749_ _1380_ net919 _1379_ VPWR VGND sg13g2_nand2_1
XFILLER_2_714 VPWR VGND sg13g2_decap_8
XFILLER_49_217 VPWR VGND sg13g2_fill_2
XFILLER_18_604 VPWR VGND sg13g2_decap_8
XFILLER_46_957 VPWR VGND sg13g2_decap_8
XFILLER_17_136 VPWR VGND sg13g2_decap_8
XFILLER_17_147 VPWR VGND sg13g2_fill_2
XFILLER_14_832 VPWR VGND sg13g2_decap_4
XFILLER_26_681 VPWR VGND sg13g2_decap_8
XFILLER_40_150 VPWR VGND sg13g2_fill_2
XFILLER_5_563 VPWR VGND sg13g2_fill_2
Xoutput1 net1 uio_out[2] VPWR VGND sg13g2_buf_1
XFILLER_49_751 VPWR VGND sg13g2_decap_8
X_4080_ net312 net1208 _2441_ VPWR VGND sg13g2_nor2_1
XFILLER_48_294 VPWR VGND sg13g2_decap_4
XFILLER_37_957 VPWR VGND sg13g2_decap_8
XFILLER_36_456 VPWR VGND sg13g2_decap_8
X_4982_ net1139 VPWR _0690_ VGND _0688_ _0689_ sg13g2_o21ai_1
XFILLER_23_128 VPWR VGND sg13g2_decap_4
XFILLER_16_191 VPWR VGND sg13g2_decap_8
X_3933_ VPWR _0252_ net459 VGND sg13g2_inv_1
X_3864_ _2198_ _2248_ _2249_ VPWR VGND sg13g2_and2_1
XFILLER_20_846 VPWR VGND sg13g2_decap_8
X_5603_ VGND VPWR _1181_ _1253_ _1254_ net1078 sg13g2_a21oi_1
X_3795_ net961 VPWR _2187_ VGND _2185_ _2186_ sg13g2_o21ai_1
X_5534_ _1191_ net1090 _1190_ VPWR VGND sg13g2_nand2b_1
X_5465_ _1126_ _1129_ net1335 _1130_ VPWR VGND sg13g2_nand3_1
X_4416_ VGND VPWR net926 _2624_ _2742_ _2741_ sg13g2_a21oi_1
XFILLER_28_1000 VPWR VGND sg13g2_decap_8
X_5396_ VGND VPWR net1103 _1064_ _1065_ _1021_ sg13g2_a21oi_1
X_4347_ net1182 net1049 _2677_ VPWR VGND sg13g2_nor2b_1
X_4278_ _2610_ VPWR _2618_ VGND _2606_ _2613_ sg13g2_o21ai_1
X_3229_ s0.data_out\[7\]\[5\] s0.data_out\[6\]\[5\] net1010 _1674_ VPWR VGND sg13g2_mux2_1
X_6017_ net267 VGND VPWR _0067_ s0.data_out\[16\]\[4\] clknet_leaf_32_clk sg13g2_dfrbpq_2
XFILLER_43_905 VPWR VGND sg13g2_decap_8
XFILLER_28_979 VPWR VGND sg13g2_decap_8
XFILLER_14_106 VPWR VGND sg13g2_decap_4
XFILLER_22_150 VPWR VGND sg13g2_decap_4
XFILLER_11_857 VPWR VGND sg13g2_decap_4
XFILLER_7_817 VPWR VGND sg13g2_decap_8
XFILLER_11_868 VPWR VGND sg13g2_fill_1
XFILLER_2_577 VPWR VGND sg13g2_decap_4
X_6019__265 VPWR VGND net265 sg13g2_tiehi
XFILLER_46_754 VPWR VGND sg13g2_decap_8
X_6165__107 VPWR VGND net107 sg13g2_tiehi
XFILLER_34_949 VPWR VGND sg13g2_decap_8
XFILLER_42_971 VPWR VGND sg13g2_decap_8
XFILLER_14_651 VPWR VGND sg13g2_fill_2
XFILLER_41_481 VPWR VGND sg13g2_fill_2
XFILLER_9_143 VPWR VGND sg13g2_decap_8
X_3580_ VGND VPWR _1991_ net511 net1313 sg13g2_or2_1
X_5250_ VGND VPWR net1107 net588 _0933_ _0932_ sg13g2_a21oi_1
X_4201_ net359 net1207 _2545_ VPWR VGND sg13g2_nor2b_1
X_5181_ _0857_ _0873_ _0874_ VPWR VGND sg13g2_nor2b_1
X_4132_ VPWR _2491_ s0.data_out\[7\]\[2\] VGND sg13g2_inv_1
X_4063_ _2424_ VPWR _2425_ VGND _2465_ net1045 sg13g2_o21ai_1
XFILLER_37_743 VPWR VGND sg13g2_decap_4
XFILLER_3_1013 VPWR VGND sg13g2_decap_8
X_4965_ VGND VPWR net1124 net386 _0675_ _0674_ sg13g2_a21oi_1
X_3916_ _2296_ VPWR _2297_ VGND net1293 net448 sg13g2_o21ai_1
X_4896_ VGND VPWR net1148 _0612_ _0613_ _0585_ sg13g2_a21oi_1
XFILLER_22_49 VPWR VGND sg13g2_fill_1
X_3847_ s0.data_out\[2\]\[2\] s0.data_out\[1\]\[2\] net955 _2232_ VPWR VGND sg13g2_mux2_1
X_3778_ _2172_ VPWR _2173_ VGND net953 _2166_ sg13g2_o21ai_1
XFILLER_4_809 VPWR VGND sg13g2_decap_8
X_5517_ VGND VPWR _1083_ _1174_ _1175_ net1093 sg13g2_a21oi_1
X_5448_ net1093 VPWR _1115_ VGND net1229 net1080 sg13g2_o21ai_1
Xfanout1109 s0.valid_out\[12\][0] net1109 VPWR VGND sg13g2_buf_1
X_5379_ net1091 net1051 _1050_ VPWR VGND sg13g2_nor2b_1
XFILLER_16_916 VPWR VGND sg13g2_fill_2
XFILLER_27_275 VPWR VGND sg13g2_decap_8
XFILLER_42_234 VPWR VGND sg13g2_fill_1
XFILLER_30_429 VPWR VGND sg13g2_fill_2
XFILLER_11_610 VPWR VGND sg13g2_fill_1
XFILLER_24_993 VPWR VGND sg13g2_decap_8
XFILLER_7_625 VPWR VGND sg13g2_decap_4
XFILLER_6_102 VPWR VGND sg13g2_fill_2
XFILLER_3_831 VPWR VGND sg13g2_decap_8
XFILLER_2_396 VPWR VGND sg13g2_fill_1
X_6032__251 VPWR VGND net251 sg13g2_tiehi
XFILLER_34_702 VPWR VGND sg13g2_fill_1
XFILLER_33_245 VPWR VGND sg13g2_fill_1
XFILLER_42_790 VPWR VGND sg13g2_fill_2
X_4750_ VGND VPWR net1160 _0478_ _0479_ _0436_ sg13g2_a21oi_1
XFILLER_21_429 VPWR VGND sg13g2_fill_2
X_3701_ VGND VPWR _2101_ net355 net1310 sg13g2_or2_1
X_4681_ net1306 VPWR _0420_ VGND net375 _0419_ sg13g2_o21ai_1
X_3632_ VGND VPWR _2041_ _2040_ net1215 sg13g2_or2_1
X_5302_ _0983_ net1111 net501 VPWR VGND sg13g2_nand2_1
X_3563_ net986 VPWR _1976_ VGND _1974_ _1975_ sg13g2_o21ai_1
XFILLER_45_0 VPWR VGND sg13g2_decap_8
X_3494_ s0.data_out\[5\]\[4\] s0.data_out\[4\]\[4\] net989 _1915_ VPWR VGND sg13g2_mux2_1
X_5233_ net1102 s0.data_out\[12\]\[4\] _0918_ VPWR VGND sg13g2_and2_1
X_5164_ _0855_ _0856_ _0854_ _0857_ VPWR VGND sg13g2_nand3_1
X_4115_ _2474_ net1239 VPWR VGND sg13g2_inv_2
X_5095_ _0793_ net937 _0792_ VPWR VGND sg13g2_nand2_1
X_4046_ VGND VPWR net941 net1061 _2412_ _2411_ sg13g2_a21oi_1
XFILLER_25_768 VPWR VGND sg13g2_decap_8
X_5997_ net289 VGND VPWR _0047_ s0.shift_out\[18\][0] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_24_278 VPWR VGND sg13g2_fill_1
X_4948_ net1122 s0.data_out\[14\]\[1\] _0660_ VPWR VGND sg13g2_and2_1
XFILLER_33_48 VPWR VGND sg13g2_fill_2
X_4879_ _0596_ net1149 _0595_ VPWR VGND sg13g2_nand2b_1
XFILLER_20_451 VPWR VGND sg13g2_fill_1
XFILLER_4_606 VPWR VGND sg13g2_decap_8
XFILLER_20_495 VPWR VGND sg13g2_decap_8
XFILLER_4_639 VPWR VGND sg13g2_fill_1
XFILLER_0_845 VPWR VGND sg13g2_decap_8
X_6016__268 VPWR VGND net268 sg13g2_tiehi
XFILLER_43_532 VPWR VGND sg13g2_decap_4
XFILLER_43_565 VPWR VGND sg13g2_fill_2
XFILLER_15_267 VPWR VGND sg13g2_decap_8
X_6199__70 VPWR VGND net70 sg13g2_tiehi
XFILLER_12_985 VPWR VGND sg13g2_decap_8
XFILLER_8_978 VPWR VGND sg13g2_decap_8
XFILLER_48_1025 VPWR VGND sg13g2_decap_4
XFILLER_39_816 VPWR VGND sg13g2_fill_1
XFILLER_47_871 VPWR VGND sg13g2_decap_8
XFILLER_0_30 VPWR VGND sg13g2_fill_1
XFILLER_0_1027 VPWR VGND sg13g2_fill_2
X_5920_ _1533_ net1013 _1493_ _1534_ VPWR VGND sg13g2_a21o_1
X_5851_ _1473_ _1474_ _1475_ VPWR VGND sg13g2_nor2b_1
X_5782_ net1027 net1047 _1409_ VPWR VGND sg13g2_nor2b_1
X_4802_ _0527_ _0528_ _0529_ VPWR VGND sg13g2_nor2_1
XFILLER_34_598 VPWR VGND sg13g2_decap_8
X_4733_ VGND VPWR _0385_ _0463_ _0464_ net1161 sg13g2_a21oi_1
X_4664_ _0392_ _0398_ _0404_ _0405_ VPWR VGND sg13g2_nor3_1
X_3615_ _2024_ net977 net576 VPWR VGND sg13g2_nand2_1
X_4595_ _0339_ s0.data_out\[17\]\[5\] net1177 VPWR VGND sg13g2_nand2b_1
X_3546_ VGND VPWR net969 net420 _1961_ _1960_ sg13g2_a21oi_1
X_5216_ _0903_ net935 _0902_ VPWR VGND sg13g2_nand2_1
X_3477_ VGND VPWR net982 _1897_ _1898_ _1851_ sg13g2_a21oi_1
X_6196_ net74 VGND VPWR _0246_ s0.shift_out\[2\][0] clknet_leaf_11_clk sg13g2_dfrbpq_2
X_5147_ _0840_ net1120 net507 VPWR VGND sg13g2_nand2_1
XFILLER_28_15 VPWR VGND sg13g2_decap_4
XFILLER_29_304 VPWR VGND sg13g2_fill_2
X_5078_ _0778_ net471 net1131 VPWR VGND sg13g2_nand2b_1
X_4029_ net1225 _2398_ _0261_ VPWR VGND sg13g2_nor2_1
XFILLER_38_882 VPWR VGND sg13g2_fill_1
XFILLER_37_392 VPWR VGND sg13g2_decap_4
XFILLER_25_587 VPWR VGND sg13g2_decap_8
XFILLER_40_546 VPWR VGND sg13g2_fill_1
XFILLER_21_793 VPWR VGND sg13g2_fill_2
XFILLER_5_937 VPWR VGND sg13g2_decap_8
XFILLER_0_642 VPWR VGND sg13g2_decap_8
XFILLER_48_668 VPWR VGND sg13g2_decap_8
XFILLER_36_808 VPWR VGND sg13g2_decap_8
XFILLER_47_189 VPWR VGND sg13g2_fill_2
XFILLER_16_543 VPWR VGND sg13g2_decap_8
XFILLER_44_885 VPWR VGND sg13g2_decap_8
XFILLER_43_395 VPWR VGND sg13g2_fill_1
XFILLER_16_598 VPWR VGND sg13g2_decap_8
XFILLER_8_753 VPWR VGND sg13g2_fill_2
XFILLER_8_775 VPWR VGND sg13g2_decap_4
Xhold208 s0.data_out\[12\]\[2\] VPWR VGND net504 sg13g2_dlygate4sd3_1
Xhold219 s0.data_out\[3\]\[7\] VPWR VGND net515 sg13g2_dlygate4sd3_1
X_4380_ _2707_ VPWR _2708_ VGND _2701_ _2702_ sg13g2_o21ai_1
X_3400_ net981 s0.data_out\[4\]\[0\] _1829_ VPWR VGND sg13g2_and2_1
X_3331_ net1325 VPWR _1765_ VGND net916 _1764_ sg13g2_o21ai_1
XFILLER_4_970 VPWR VGND sg13g2_decap_8
X_3262_ VPWR _1705_ _1704_ VGND sg13g2_inv_1
X_6050_ net231 VGND VPWR _0100_ s0.data_out\[13\]\[1\] clknet_leaf_29_clk sg13g2_dfrbpq_2
X_3193_ net1326 VPWR _1640_ VGND net917 _1639_ sg13g2_o21ai_1
XFILLER_39_635 VPWR VGND sg13g2_fill_1
X_5001_ VPWR _0082_ net555 VGND sg13g2_inv_1
XFILLER_22_1006 VPWR VGND sg13g2_decap_8
XFILLER_38_123 VPWR VGND sg13g2_fill_1
Xfanout1270 net1271 net1270 VPWR VGND sg13g2_buf_8
Xfanout1281 net1284 net1281 VPWR VGND sg13g2_buf_8
Xfanout1292 net1296 net1292 VPWR VGND sg13g2_buf_8
XFILLER_26_318 VPWR VGND sg13g2_fill_2
XFILLER_38_189 VPWR VGND sg13g2_fill_2
X_5903_ _1519_ net544 net1032 VPWR VGND sg13g2_nand2b_1
X_5834_ VGND VPWR _1394_ _1453_ _1460_ net1252 sg13g2_a21oi_1
XFILLER_34_373 VPWR VGND sg13g2_decap_8
X_5765_ _1394_ net920 _1393_ VPWR VGND sg13g2_nand2_1
X_4716_ s0.data_out\[16\]\[4\] s0.data_out\[17\]\[4\] net1165 _0449_ VPWR VGND sg13g2_mux2_1
X_5696_ _1327_ _1340_ _1313_ _1341_ VPWR VGND sg13g2_nand3_1
X_4647_ VGND VPWR net1171 _0387_ _0388_ _0347_ sg13g2_a21oi_1
X_4578_ VPWR _0041_ net499 VGND sg13g2_inv_1
X_3529_ net969 s0.data_out\[3\]\[0\] _1946_ VPWR VGND sg13g2_and2_1
X_6179_ net92 VGND VPWR _0229_ s0.data_out\[3\]\[3\] clknet_leaf_6_clk sg13g2_dfrbpq_2
XFILLER_38_690 VPWR VGND sg13g2_decap_4
XFILLER_26_852 VPWR VGND sg13g2_decap_8
XFILLER_26_863 VPWR VGND sg13g2_fill_2
XFILLER_41_822 VPWR VGND sg13g2_decap_8
XFILLER_38_1024 VPWR VGND sg13g2_decap_4
XFILLER_13_535 VPWR VGND sg13g2_decap_4
XFILLER_25_362 VPWR VGND sg13g2_decap_4
XFILLER_25_384 VPWR VGND sg13g2_fill_2
XFILLER_26_885 VPWR VGND sg13g2_decap_8
X_6184__87 VPWR VGND net87 sg13g2_tiehi
XFILLER_4_288 VPWR VGND sg13g2_decap_4
XFILLER_45_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_933 VPWR VGND sg13g2_decap_8
XFILLER_1_984 VPWR VGND sg13g2_decap_8
XFILLER_48_443 VPWR VGND sg13g2_decap_8
Xhold91 s0.data_out\[15\]\[3\] VPWR VGND net387 sg13g2_dlygate4sd3_1
Xhold80 _0049_ VPWR VGND net376 sg13g2_dlygate4sd3_1
XFILLER_35_137 VPWR VGND sg13g2_fill_2
XFILLER_32_800 VPWR VGND sg13g2_fill_1
XFILLER_44_671 VPWR VGND sg13g2_decap_4
XFILLER_32_833 VPWR VGND sg13g2_decap_4
X_3880_ s0.data_out\[2\]\[4\] s0.data_out\[1\]\[4\] net958 _2265_ VPWR VGND sg13g2_mux2_1
XFILLER_16_395 VPWR VGND sg13g2_fill_1
XFILLER_31_332 VPWR VGND sg13g2_decap_4
XFILLER_31_376 VPWR VGND sg13g2_fill_2
XFILLER_12_590 VPWR VGND sg13g2_fill_2
X_5550_ _1207_ _1206_ net1242 _1202_ net1236 VPWR VGND sg13g2_a22oi_1
X_4501_ net1284 _2816_ _2817_ VPWR VGND sg13g2_nor2b_1
X_5481_ VGND VPWR _1144_ net568 net1337 sg13g2_or2_1
X_4432_ _2693_ VPWR _2755_ VGND net1187 _2484_ sg13g2_o21ai_1
X_4363_ VGND VPWR net1193 _2690_ _2691_ _2648_ sg13g2_a21oi_1
XFILLER_6_95 VPWR VGND sg13g2_decap_8
X_3314_ VGND VPWR net995 net352 _1750_ _1749_ sg13g2_a21oi_1
X_6102_ net176 VGND VPWR _0152_ s0.was_valid_out\[9\][0] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_4294_ net1289 VPWR _2632_ VGND net435 _2626_ sg13g2_o21ai_1
X_3245_ VGND VPWR net1015 _1689_ _1690_ _1637_ sg13g2_a21oi_1
X_6033_ net250 VGND VPWR _0083_ s0.shift_out\[15\][0] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_3176_ VGND VPWR net1005 net423 _1625_ _1624_ sg13g2_a21oi_1
XFILLER_39_498 VPWR VGND sg13g2_fill_1
XFILLER_41_118 VPWR VGND sg13g2_fill_1
XFILLER_22_310 VPWR VGND sg13g2_fill_1
X_5817_ VGND VPWR net1037 _1442_ _1443_ _1401_ sg13g2_a21oi_1
X_5748_ s0.data_out\[8\]\[3\] s0.data_out\[9\]\[3\] net1041 _1379_ VPWR VGND sg13g2_mux2_1
X_5679_ net1243 _1321_ _1324_ VPWR VGND sg13g2_nor2_1
XFILLER_46_936 VPWR VGND sg13g2_decap_8
XFILLER_13_321 VPWR VGND sg13g2_fill_1
XFILLER_41_685 VPWR VGND sg13g2_fill_1
XFILLER_41_663 VPWR VGND sg13g2_fill_2
XFILLER_40_162 VPWR VGND sg13g2_decap_8
XFILLER_13_354 VPWR VGND sg13g2_decap_8
XFILLER_13_365 VPWR VGND sg13g2_fill_2
XFILLER_15_93 VPWR VGND sg13g2_fill_2
XFILLER_12_1027 VPWR VGND sg13g2_fill_2
XFILLER_49_7 VPWR VGND sg13g2_decap_8
Xoutput2 net2 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_1_781 VPWR VGND sg13g2_decap_8
XFILLER_49_730 VPWR VGND sg13g2_decap_8
XFILLER_37_936 VPWR VGND sg13g2_decap_8
XFILLER_36_435 VPWR VGND sg13g2_decap_8
XFILLER_45_991 VPWR VGND sg13g2_decap_8
X_4981_ net1125 net1055 _0689_ VPWR VGND sg13g2_nor2b_1
X_3932_ _2310_ VPWR _2311_ VGND net1293 net458 sg13g2_o21ai_1
X_3863_ _2248_ net961 _2247_ VPWR VGND sg13g2_nand2b_1
X_5602_ _1253_ net451 net1084 VPWR VGND sg13g2_nand2b_1
X_5533_ VGND VPWR net1077 _1189_ _1190_ _1128_ sg13g2_a21oi_1
X_3794_ net949 net1069 _2186_ VPWR VGND sg13g2_nor2b_1
XFILLER_8_391 VPWR VGND sg13g2_decap_4
X_5464_ net1090 VPWR _1129_ VGND _1127_ _1128_ sg13g2_o21ai_1
X_4415_ _2739_ _2740_ _2741_ VPWR VGND sg13g2_nor2_1
X_5395_ _1063_ net1089 _1022_ _1064_ VPWR VGND sg13g2_a21o_1
X_4346_ VGND VPWR _2595_ _2675_ _2676_ net1197 sg13g2_a21oi_1
X_4277_ _2599_ _2600_ _2617_ VPWR VGND sg13g2_nor2_1
X_3228_ _1673_ net1009 net539 VPWR VGND sg13g2_nand2_1
XFILLER_39_240 VPWR VGND sg13g2_fill_2
X_6016_ net268 VGND VPWR _0066_ s0.data_out\[16\]\[3\] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_3159_ net1001 s0.data_out\[6\]\[2\] _1610_ VPWR VGND sg13g2_and2_1
XFILLER_28_969 VPWR VGND sg13g2_fill_1
XFILLER_36_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_34_clk clknet_3_1__leaf_clk clknet_leaf_34_clk VPWR VGND sg13g2_buf_8
XFILLER_35_1027 VPWR VGND sg13g2_fill_2
XFILLER_11_803 VPWR VGND sg13g2_decap_8
XFILLER_11_814 VPWR VGND sg13g2_fill_2
XFILLER_7_807 VPWR VGND sg13g2_fill_1
XFILLER_10_302 VPWR VGND sg13g2_decap_8
X_6158__115 VPWR VGND net115 sg13g2_tiehi
XFILLER_2_556 VPWR VGND sg13g2_decap_8
XFILLER_46_733 VPWR VGND sg13g2_decap_8
XFILLER_18_402 VPWR VGND sg13g2_decap_8
XFILLER_45_243 VPWR VGND sg13g2_decap_8
XFILLER_34_906 VPWR VGND sg13g2_fill_2
XFILLER_45_276 VPWR VGND sg13g2_decap_8
XFILLER_42_950 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_25_clk clknet_3_5__leaf_clk clknet_leaf_25_clk VPWR VGND sg13g2_buf_8
XFILLER_33_438 VPWR VGND sg13g2_decap_4
XFILLER_14_685 VPWR VGND sg13g2_decap_8
XFILLER_9_199 VPWR VGND sg13g2_fill_2
XFILLER_10_880 VPWR VGND sg13g2_fill_1
XFILLER_6_884 VPWR VGND sg13g2_decap_8
X_4200_ net1204 VPWR _2544_ VGND _2542_ _2543_ sg13g2_o21ai_1
X_5180_ _0870_ VPWR _0873_ VGND _0861_ _0866_ sg13g2_o21ai_1
X_4131_ _2490_ s0.data_out\[9\]\[5\] VPWR VGND sg13g2_inv_2
X_4062_ net334 net947 net944 _2424_ VPWR VGND sg13g2_a21o_1
XFILLER_18_980 VPWR VGND sg13g2_decap_8
XFILLER_40_909 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_16_clk clknet_3_6__leaf_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
X_4964_ net1124 net1063 _0674_ VPWR VGND sg13g2_nor2b_1
X_3915_ _2292_ _2295_ net1293 _2296_ VPWR VGND sg13g2_nand3_1
XFILLER_33_983 VPWR VGND sg13g2_decap_8
X_4895_ _0611_ net1136 _0586_ _0612_ VPWR VGND sg13g2_a21o_1
X_3846_ VPWR _0245_ _2231_ VGND sg13g2_inv_1
XFILLER_20_666 VPWR VGND sg13g2_decap_4
X_3777_ net930 VPWR _2172_ VGND net328 net966 sg13g2_o21ai_1
X_5516_ _1174_ net531 net1097 VPWR VGND sg13g2_nand2b_1
X_5447_ net316 net1345 _0120_ VPWR VGND sg13g2_and2_1
X_5378_ VGND VPWR _0969_ _1048_ _1049_ net1105 sg13g2_a21oi_1
X_4329_ s0.data_out\[19\]\[4\] s0.data_out\[20\]\[4\] net1200 _2661_ VPWR VGND sg13g2_mux2_1
XFILLER_47_14 VPWR VGND sg13g2_decap_8
XFILLER_27_221 VPWR VGND sg13g2_fill_1
XFILLER_24_972 VPWR VGND sg13g2_decap_8
XFILLER_10_143 VPWR VGND sg13g2_decap_4
XFILLER_11_688 VPWR VGND sg13g2_fill_2
XFILLER_12_61 VPWR VGND sg13g2_fill_2
XFILLER_3_810 VPWR VGND sg13g2_decap_8
X_6171__101 VPWR VGND net101 sg13g2_tiehi
XFILLER_3_887 VPWR VGND sg13g2_decap_8
XFILLER_33_202 VPWR VGND sg13g2_decap_8
XFILLER_34_714 VPWR VGND sg13g2_fill_1
XFILLER_34_747 VPWR VGND sg13g2_fill_2
XFILLER_18_1022 VPWR VGND sg13g2_decap_8
XFILLER_21_419 VPWR VGND sg13g2_fill_2
X_3700_ net1309 VPWR _2100_ VGND net933 _2099_ sg13g2_o21ai_1
XFILLER_15_994 VPWR VGND sg13g2_decap_8
X_4680_ _0414_ VPWR _0419_ VGND net1159 _0295_ sg13g2_o21ai_1
X_3631_ _1973_ VPWR _2040_ VGND net914 _2039_ sg13g2_o21ai_1
X_3562_ net970 net1058 _1975_ VPWR VGND sg13g2_nor2b_1
X_5301_ VGND VPWR _0982_ _0981_ net1215 sg13g2_or2_1
X_3493_ _1912_ _1913_ _1911_ _1914_ VPWR VGND sg13g2_nand3_1
X_5232_ _0917_ net935 _0916_ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_5_clk clknet_3_6__leaf_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
XFILLER_38_0 VPWR VGND sg13g2_decap_8
X_5163_ VGND VPWR _0856_ _0853_ net1242 sg13g2_or2_1
X_4114_ VPWR _2473_ net356 VGND sg13g2_inv_1
X_5094_ s0.data_out\[13\]\[3\] s0.data_out\[14\]\[3\] net1131 _0792_ VPWR VGND sg13g2_mux2_1
X_4045_ net941 _2361_ _2411_ VPWR VGND sg13g2_nor2_1
XFILLER_25_747 VPWR VGND sg13g2_decap_8
X_5996_ net290 VGND VPWR _0046_ s0.data_out\[18\]\[7\] clknet_leaf_35_clk sg13g2_dfrbpq_2
XFILLER_40_739 VPWR VGND sg13g2_fill_1
X_4947_ _0659_ net921 _0658_ VPWR VGND sg13g2_nand2_1
XFILLER_21_920 VPWR VGND sg13g2_decap_8
X_4878_ VGND VPWR net1135 _0594_ _0595_ _0545_ sg13g2_a21oi_1
X_6009__276 VPWR VGND net276 sg13g2_tiehi
X_3829_ _2216_ VPWR _2217_ VGND net1299 net349 sg13g2_o21ai_1
XFILLER_20_485 VPWR VGND sg13g2_fill_1
XFILLER_21_997 VPWR VGND sg13g2_decap_8
XFILLER_3_106 VPWR VGND sg13g2_fill_2
X_6155__118 VPWR VGND net118 sg13g2_tiehi
XFILLER_0_824 VPWR VGND sg13g2_decap_8
XFILLER_15_246 VPWR VGND sg13g2_decap_8
XFILLER_31_739 VPWR VGND sg13g2_decap_8
XFILLER_12_964 VPWR VGND sg13g2_decap_8
XFILLER_8_957 VPWR VGND sg13g2_decap_8
XFILLER_48_1004 VPWR VGND sg13g2_decap_8
XFILLER_39_839 VPWR VGND sg13g2_fill_2
XFILLER_38_305 VPWR VGND sg13g2_fill_2
XFILLER_47_850 VPWR VGND sg13g2_decap_8
XFILLER_19_530 VPWR VGND sg13g2_fill_2
XFILLER_0_1006 VPWR VGND sg13g2_decap_8
X_5850_ net918 VPWR _1474_ VGND net326 net1032 sg13g2_o21ai_1
XFILLER_0_97 VPWR VGND sg13g2_fill_2
X_5781_ VGND VPWR _1314_ _1407_ _1408_ net1038 sg13g2_a21oi_1
X_4801_ VGND VPWR net1222 net1153 _0528_ net1148 sg13g2_a21oi_1
XFILLER_22_739 VPWR VGND sg13g2_decap_8
X_4732_ _0463_ net546 net1165 VPWR VGND sg13g2_nand2b_1
X_4663_ net1248 _0396_ _0404_ VPWR VGND sg13g2_nor2_1
XFILLER_30_761 VPWR VGND sg13g2_decap_8
X_3614_ VGND VPWR net983 _2022_ _2023_ _1994_ sg13g2_a21oi_1
X_4594_ VPWR _0043_ _0338_ VGND sg13g2_inv_1
X_3545_ net969 net1068 _1960_ VPWR VGND sg13g2_nor2b_1
X_3476_ s0.data_out\[5\]\[3\] s0.data_out\[4\]\[3\] net989 _1897_ VPWR VGND sg13g2_mux2_1
X_5215_ s0.data_out\[12\]\[2\] s0.data_out\[13\]\[2\] net1121 _0902_ VPWR VGND sg13g2_mux2_1
XFILLER_9_1020 VPWR VGND sg13g2_decap_8
X_6195_ net75 VGND VPWR _0245_ s0.data_out\[2\]\[7\] clknet_leaf_10_clk sg13g2_dfrbpq_2
X_5146_ _0830_ _0837_ _0838_ _0839_ VPWR VGND sg13g2_nor3_1
XFILLER_45_809 VPWR VGND sg13g2_decap_8
XFILLER_38_850 VPWR VGND sg13g2_fill_2
X_5077_ VPWR _0087_ _0777_ VGND sg13g2_inv_1
X_4028_ _2397_ _2398_ _0260_ VPWR VGND sg13g2_nor2_1
XFILLER_44_319 VPWR VGND sg13g2_decap_4
X_5979_ net36 VGND VPWR _0029_ s0.data_out\[19\]\[2\] clknet_leaf_36_clk sg13g2_dfrbpq_2
XFILLER_12_205 VPWR VGND sg13g2_decap_4
X_6196__74 VPWR VGND net74 sg13g2_tiehi
XFILLER_5_916 VPWR VGND sg13g2_decap_8
X_6022__262 VPWR VGND net262 sg13g2_tiehi
XFILLER_0_621 VPWR VGND sg13g2_decap_8
XFILLER_0_698 VPWR VGND sg13g2_decap_8
XFILLER_48_647 VPWR VGND sg13g2_decap_8
XFILLER_47_179 VPWR VGND sg13g2_fill_1
XFILLER_44_864 VPWR VGND sg13g2_decap_8
XFILLER_43_385 VPWR VGND sg13g2_fill_1
XFILLER_43_374 VPWR VGND sg13g2_decap_4
XFILLER_12_761 VPWR VGND sg13g2_fill_2
XFILLER_11_293 VPWR VGND sg13g2_decap_4
XFILLER_7_242 VPWR VGND sg13g2_fill_2
Xhold209 _1026_ VPWR VGND net505 sg13g2_dlygate4sd3_1
X_3330_ VGND VPWR net995 s0.data_out\[5\]\[7\] _1764_ _1763_ sg13g2_a21oi_1
X_3261_ _1702_ _1703_ _1704_ VPWR VGND sg13g2_nor2_1
XFILLER_3_492 VPWR VGND sg13g2_fill_1
X_5000_ _0705_ VPWR _0706_ VGND _0701_ _0704_ sg13g2_o21ai_1
X_3192_ VGND VPWR net1006 s0.data_out\[6\]\[6\] _1639_ _1638_ sg13g2_a21oi_1
Xfanout1282 net1284 net1282 VPWR VGND sg13g2_buf_8
Xfanout1271 net1272 net1271 VPWR VGND sg13g2_buf_8
Xfanout1260 net1263 net1260 VPWR VGND sg13g2_buf_8
XFILLER_38_179 VPWR VGND sg13g2_fill_1
Xfanout1293 net1296 net1293 VPWR VGND sg13g2_buf_8
XFILLER_35_842 VPWR VGND sg13g2_decap_8
XFILLER_19_382 VPWR VGND sg13g2_fill_2
X_5902_ VPWR _0171_ net483 VGND sg13g2_inv_1
X_5833_ _1454_ _1458_ _1459_ VPWR VGND sg13g2_and2_1
XFILLER_22_514 VPWR VGND sg13g2_decap_8
X_5764_ s0.data_out\[8\]\[5\] s0.data_out\[9\]\[5\] net1042 _1393_ VPWR VGND sg13g2_mux2_1
X_4715_ VPWR _0054_ _0448_ VGND sg13g2_inv_1
X_5695_ _1336_ _1337_ _1338_ _1339_ _1340_ VPWR VGND sg13g2_nor4_1
X_4646_ _0386_ net1158 _0348_ _0387_ VPWR VGND sg13g2_a21o_1
X_6006__279 VPWR VGND net279 sg13g2_tiehi
XFILLER_30_28 VPWR VGND sg13g2_decap_4
X_6193__77 VPWR VGND net77 sg13g2_tiehi
X_4577_ _0323_ VPWR _0324_ VGND _0319_ _0322_ sg13g2_o21ai_1
XFILLER_1_429 VPWR VGND sg13g2_decap_8
X_3528_ _1945_ net914 _1944_ VPWR VGND sg13g2_nand2_1
X_3459_ VGND VPWR _1881_ net569 net1314 sg13g2_or2_1
X_6178_ net93 VGND VPWR _0228_ s0.data_out\[3\]\[2\] clknet_leaf_6_clk sg13g2_dfrbpq_2
X_5129_ VGND VPWR net1112 s0.data_out\[13\]\[7\] _0823_ _0822_ sg13g2_a21oi_1
XFILLER_29_168 VPWR VGND sg13g2_fill_1
XFILLER_44_127 VPWR VGND sg13g2_fill_1
XFILLER_38_1003 VPWR VGND sg13g2_decap_8
XFILLER_20_72 VPWR VGND sg13g2_fill_1
X_6096__182 VPWR VGND net182 sg13g2_tiehi
XFILLER_1_963 VPWR VGND sg13g2_decap_8
XFILLER_49_912 VPWR VGND sg13g2_decap_8
XFILLER_0_473 VPWR VGND sg13g2_fill_1
XFILLER_48_422 VPWR VGND sg13g2_decap_8
XFILLER_49_989 VPWR VGND sg13g2_decap_8
XFILLER_36_628 VPWR VGND sg13g2_decap_8
Xhold70 s0.data_out\[21\]\[3\] VPWR VGND net366 sg13g2_dlygate4sd3_1
Xhold92 s0.data_out\[21\]\[2\] VPWR VGND net388 sg13g2_dlygate4sd3_1
Xhold81 s0.data_out\[0\]\[0\] VPWR VGND net377 sg13g2_dlygate4sd3_1
XFILLER_48_499 VPWR VGND sg13g2_decap_8
XFILLER_45_91 VPWR VGND sg13g2_fill_2
XFILLER_8_573 VPWR VGND sg13g2_decap_8
X_4500_ _2749_ VPWR _2816_ VGND net926 _2815_ sg13g2_o21ai_1
X_5480_ net1344 VPWR _1143_ VGND net939 _1142_ sg13g2_o21ai_1
XFILLER_8_595 VPWR VGND sg13g2_fill_2
X_4431_ VPWR _0027_ _2754_ VGND sg13g2_inv_1
X_4362_ _2689_ net1178 _2649_ _2690_ VPWR VGND sg13g2_a21o_1
X_3313_ net995 net1055 _1749_ VPWR VGND sg13g2_nor2b_1
X_4293_ _2629_ _2630_ _2631_ VPWR VGND sg13g2_nor2b_1
X_6101_ net177 VGND VPWR _0151_ s0.data_new_delayed\[7\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_3244_ _1688_ net1006 _1638_ _1689_ VPWR VGND sg13g2_a21o_1
XFILLER_39_411 VPWR VGND sg13g2_fill_1
X_6032_ net251 VGND VPWR _0082_ s0.data_out\[15\]\[7\] clknet_leaf_30_clk sg13g2_dfrbpq_2
X_3175_ net1005 net1059 _1624_ VPWR VGND sg13g2_nor2b_1
Xfanout1090 net1095 net1090 VPWR VGND sg13g2_buf_8
XFILLER_27_606 VPWR VGND sg13g2_fill_1
X_6012__272 VPWR VGND net272 sg13g2_tiehi
XFILLER_25_39 VPWR VGND sg13g2_fill_1
XFILLER_23_856 VPWR VGND sg13g2_fill_1
X_5816_ _1441_ net1028 _1402_ _1442_ VPWR VGND sg13g2_a21o_1
XFILLER_22_377 VPWR VGND sg13g2_fill_1
XFILLER_23_878 VPWR VGND sg13g2_fill_2
XFILLER_10_528 VPWR VGND sg13g2_fill_1
X_5747_ VPWR _0156_ _1378_ VGND sg13g2_inv_1
X_5678_ VPWR _1323_ _1322_ VGND sg13g2_inv_1
X_4629_ VGND VPWR net1155 _0369_ _0370_ _0307_ sg13g2_a21oi_1
XFILLER_2_749 VPWR VGND sg13g2_decap_8
XFILLER_49_219 VPWR VGND sg13g2_fill_1
XFILLER_46_915 VPWR VGND sg13g2_decap_8
XFILLER_45_458 VPWR VGND sg13g2_fill_1
XFILLER_41_620 VPWR VGND sg13g2_decap_8
XFILLER_15_50 VPWR VGND sg13g2_fill_1
XFILLER_25_182 VPWR VGND sg13g2_fill_2
XFILLER_26_694 VPWR VGND sg13g2_fill_1
XFILLER_40_152 VPWR VGND sg13g2_fill_1
XFILLER_9_304 VPWR VGND sg13g2_decap_8
XFILLER_12_1006 VPWR VGND sg13g2_decap_8
XFILLER_31_71 VPWR VGND sg13g2_fill_1
XFILLER_5_565 VPWR VGND sg13g2_fill_1
XFILLER_31_82 VPWR VGND sg13g2_fill_2
Xoutput3 net3 uo_out[1] VPWR VGND sg13g2_buf_1
X_6180__91 VPWR VGND net91 sg13g2_tiehi
XFILLER_1_760 VPWR VGND sg13g2_decap_8
XFILLER_49_786 VPWR VGND sg13g2_decap_8
XFILLER_37_926 VPWR VGND sg13g2_fill_1
XFILLER_45_970 VPWR VGND sg13g2_decap_8
XFILLER_17_672 VPWR VGND sg13g2_fill_2
X_4980_ net1125 s0.data_out\[14\]\[5\] _0688_ VPWR VGND sg13g2_and2_1
XFILLER_23_108 VPWR VGND sg13g2_decap_8
XFILLER_16_182 VPWR VGND sg13g2_decap_4
X_3931_ _2306_ _2309_ net1292 _2310_ VPWR VGND sg13g2_nand3_1
XFILLER_31_141 VPWR VGND sg13g2_fill_1
X_3862_ VGND VPWR net950 _2246_ _2247_ _2200_ sg13g2_a21oi_1
X_5601_ VPWR _0136_ _1252_ VGND sg13g2_inv_1
X_5532_ s0.data_out\[11\]\[0\] s0.data_out\[10\]\[0\] net1084 _1189_ VPWR VGND sg13g2_mux2_1
X_3793_ net949 s0.data_out\[1\]\[1\] _2185_ VPWR VGND sg13g2_and2_1
XFILLER_9_882 VPWR VGND sg13g2_fill_1
X_5463_ net1077 net1074 _1128_ VPWR VGND sg13g2_nor2b_1
X_4414_ net1226 net1176 _2740_ VPWR VGND sg13g2_nor2b_1
X_5394_ s0.data_out\[12\]\[2\] s0.data_out\[11\]\[2\] net1096 _1063_ VPWR VGND sg13g2_mux2_1
X_4345_ _2675_ net551 net1201 VPWR VGND sg13g2_nand2b_1
X_4276_ _2590_ _2602_ _2611_ _2615_ _2616_ VPWR VGND sg13g2_or4_1
X_3227_ VGND VPWR net1015 _1671_ _1672_ _1623_ sg13g2_a21oi_1
X_6015_ net269 VGND VPWR _0065_ s0.data_out\[16\]\[2\] clknet_leaf_34_clk sg13g2_dfrbpq_2
XFILLER_28_948 VPWR VGND sg13g2_fill_1
X_3158_ _1609_ net917 _1608_ VPWR VGND sg13g2_nand2_1
XFILLER_27_447 VPWR VGND sg13g2_decap_8
XFILLER_35_1006 VPWR VGND sg13g2_decap_8
X_6086__192 VPWR VGND net192 sg13g2_tiehi
XFILLER_10_347 VPWR VGND sg13g2_fill_2
XFILLER_6_318 VPWR VGND sg13g2_decap_8
XFILLER_10_369 VPWR VGND sg13g2_fill_2
X_6093__185 VPWR VGND net185 sg13g2_tiehi
XFILLER_46_712 VPWR VGND sg13g2_decap_8
XFILLER_19_959 VPWR VGND sg13g2_decap_8
XFILLER_18_447 VPWR VGND sg13g2_decap_4
XFILLER_46_789 VPWR VGND sg13g2_decap_8
XFILLER_26_60 VPWR VGND sg13g2_fill_2
XFILLER_26_93 VPWR VGND sg13g2_decap_8
XFILLER_14_653 VPWR VGND sg13g2_fill_1
XFILLER_6_841 VPWR VGND sg13g2_decap_4
X_4130_ VPWR _2489_ s0.data_out\[9\]\[2\] VGND sg13g2_inv_1
X_4061_ net1294 net334 _2423_ VPWR VGND sg13g2_nor2_1
XFILLER_49_583 VPWR VGND sg13g2_decap_8
X_4963_ _0673_ net921 _0672_ VPWR VGND sg13g2_nand2_1
XFILLER_17_480 VPWR VGND sg13g2_fill_2
X_5959__58 VPWR VGND net58 sg13g2_tiehi
X_3914_ net951 VPWR _2295_ VGND _2293_ _2294_ sg13g2_o21ai_1
XFILLER_33_962 VPWR VGND sg13g2_decap_8
X_4894_ s0.data_out\[16\]\[7\] s0.data_out\[15\]\[7\] net1141 _0611_ VPWR VGND sg13g2_mux2_1
XFILLER_32_483 VPWR VGND sg13g2_decap_8
X_3845_ _2230_ VPWR _2231_ VGND _2226_ _2229_ sg13g2_o21ai_1
X_3776_ _2168_ VPWR _2171_ VGND net328 net957 sg13g2_o21ai_1
X_5515_ VPWR _0129_ _1173_ VGND sg13g2_inv_1
X_5446_ VGND VPWR _1109_ _1113_ _0119_ _1114_ sg13g2_a21oi_1
X_5377_ _1048_ net527 net1110 VPWR VGND sg13g2_nand2b_1
X_4328_ VPWR _0018_ net561 VGND sg13g2_inv_1
XFILLER_41_1010 VPWR VGND sg13g2_decap_8
X_4259_ _2599_ _2598_ net1239 _2594_ net1231 VPWR VGND sg13g2_a22oi_1
XFILLER_28_712 VPWR VGND sg13g2_fill_1
XFILLER_27_244 VPWR VGND sg13g2_fill_2
XFILLER_28_756 VPWR VGND sg13g2_fill_2
XFILLER_15_417 VPWR VGND sg13g2_decap_4
XFILLER_16_918 VPWR VGND sg13g2_fill_1
XFILLER_43_737 VPWR VGND sg13g2_decap_8
XFILLER_11_656 VPWR VGND sg13g2_decap_4
XFILLER_23_494 VPWR VGND sg13g2_decap_8
XFILLER_7_649 VPWR VGND sg13g2_decap_4
XFILLER_6_104 VPWR VGND sg13g2_fill_1
XFILLER_10_177 VPWR VGND sg13g2_fill_2
XFILLER_6_159 VPWR VGND sg13g2_fill_1
XFILLER_3_866 VPWR VGND sg13g2_decap_8
XFILLER_2_343 VPWR VGND sg13g2_decap_8
XFILLER_19_767 VPWR VGND sg13g2_fill_2
XFILLER_46_553 VPWR VGND sg13g2_decap_4
XFILLER_18_266 VPWR VGND sg13g2_fill_1
XFILLER_18_1001 VPWR VGND sg13g2_decap_8
XFILLER_42_792 VPWR VGND sg13g2_fill_1
XFILLER_42_770 VPWR VGND sg13g2_fill_2
XFILLER_14_483 VPWR VGND sg13g2_fill_1
XFILLER_14_494 VPWR VGND sg13g2_fill_2
X_3630_ VGND VPWR net970 _2038_ _2039_ _1975_ sg13g2_a21oi_1
X_3561_ net970 s0.data_out\[3\]\[4\] _1974_ VPWR VGND sg13g2_and2_1
X_5300_ _0917_ VPWR _0981_ VGND net935 _0980_ sg13g2_o21ai_1
X_3492_ VGND VPWR _1913_ _1910_ net1240 sg13g2_or2_1
XFILLER_5_181 VPWR VGND sg13g2_fill_1
X_5231_ s0.data_out\[12\]\[4\] s0.data_out\[13\]\[4\] net1120 _0916_ VPWR VGND sg13g2_mux2_1
X_5162_ VGND VPWR _0855_ _0849_ net1236 sg13g2_or2_1
X_5093_ VPWR _0089_ _0791_ VGND sg13g2_inv_1
X_4113_ VPWR _2472_ net364 VGND sg13g2_inv_1
XFILLER_25_1027 VPWR VGND sg13g2_fill_2
XFILLER_49_380 VPWR VGND sg13g2_decap_8
X_4044_ net1292 net348 _2410_ VPWR VGND sg13g2_nor2_1
X_6148__126 VPWR VGND net126 sg13g2_tiehi
X_5995_ net291 VGND VPWR _0045_ s0.data_out\[18\]\[6\] clknet_leaf_33_clk sg13g2_dfrbpq_2
XFILLER_24_258 VPWR VGND sg13g2_decap_8
X_4946_ s0.data_out\[14\]\[1\] s0.data_out\[15\]\[1\] net1142 _0658_ VPWR VGND sg13g2_mux2_1
X_4877_ s0.data_out\[16\]\[1\] s0.data_out\[15\]\[1\] net1141 _0594_ VPWR VGND sg13g2_mux2_1
XFILLER_21_954 VPWR VGND sg13g2_fill_1
X_3828_ _2212_ _2215_ net1299 _2216_ VPWR VGND sg13g2_nand3_1
X_3759_ net1248 _2154_ _2156_ VPWR VGND sg13g2_nor2_1
XFILLER_0_803 VPWR VGND sg13g2_decap_8
X_5429_ VGND VPWR net1103 _1097_ _1098_ _1035_ sg13g2_a21oi_1
XFILLER_48_829 VPWR VGND sg13g2_decap_8
XFILLER_47_317 VPWR VGND sg13g2_decap_4
X_6090__188 VPWR VGND net188 sg13g2_tiehi
XFILLER_16_715 VPWR VGND sg13g2_decap_8
XFILLER_15_225 VPWR VGND sg13g2_fill_2
XFILLER_16_737 VPWR VGND sg13g2_fill_1
XFILLER_28_597 VPWR VGND sg13g2_decap_8
XFILLER_31_718 VPWR VGND sg13g2_fill_1
XFILLER_43_589 VPWR VGND sg13g2_fill_2
XFILLER_12_943 VPWR VGND sg13g2_decap_8
XFILLER_8_936 VPWR VGND sg13g2_decap_8
XFILLER_11_464 VPWR VGND sg13g2_decap_4
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_19_575 VPWR VGND sg13g2_decap_8
XFILLER_34_501 VPWR VGND sg13g2_decap_8
XFILLER_34_512 VPWR VGND sg13g2_fill_2
XFILLER_34_523 VPWR VGND sg13g2_fill_1
X_4800_ _0525_ _0526_ _0527_ VPWR VGND sg13g2_nor2_2
X_5780_ _1407_ s0.data_out\[8\]\[7\] net1043 VPWR VGND sg13g2_nand2b_1
X_4731_ VPWR _0056_ net583 VGND sg13g2_inv_1
X_4662_ _0333_ _0401_ net1255 _0403_ VPWR VGND sg13g2_nand3_1
X_3613_ _2021_ net972 _1995_ _2022_ VPWR VGND sg13g2_a21o_1
XFILLER_31_1020 VPWR VGND sg13g2_decap_8
X_4593_ _0337_ VPWR _0338_ VGND net1303 net325 sg13g2_o21ai_1
X_3544_ VGND VPWR _1883_ _1958_ _1959_ net980 sg13g2_a21oi_1
X_3475_ _1887_ VPWR _1896_ VGND net1280 _1891_ sg13g2_o21ai_1
X_5214_ VPWR _0100_ _0901_ VGND sg13g2_inv_1
X_6194_ net76 VGND VPWR _0244_ s0.data_out\[2\]\[6\] clknet_leaf_10_clk sg13g2_dfrbpq_2
X_5145_ VPWR VGND _0772_ net1283 _0836_ net1279 _0838_ _0833_ sg13g2_a221oi_1
XFILLER_29_306 VPWR VGND sg13g2_fill_1
X_5076_ _0776_ VPWR _0777_ VGND net1321 net457 sg13g2_o21ai_1
X_4027_ net1294 VPWR _2398_ VGND net947 net944 sg13g2_o21ai_1
XFILLER_37_350 VPWR VGND sg13g2_decap_8
X_6161__112 VPWR VGND net112 sg13g2_tiehi
XFILLER_40_504 VPWR VGND sg13g2_decap_8
X_5978_ net37 VGND VPWR _0028_ s0.data_out\[19\]\[1\] clknet_leaf_36_clk sg13g2_dfrbpq_2
XFILLER_40_537 VPWR VGND sg13g2_fill_2
X_4929_ net1140 _0526_ _0644_ VPWR VGND sg13g2_nor2_1
XFILLER_21_784 VPWR VGND sg13g2_decap_4
XFILLER_4_438 VPWR VGND sg13g2_decap_4
XFILLER_0_600 VPWR VGND sg13g2_decap_8
XFILLER_48_626 VPWR VGND sg13g2_decap_8
XFILLER_0_677 VPWR VGND sg13g2_decap_8
XFILLER_29_862 VPWR VGND sg13g2_decap_8
XFILLER_44_843 VPWR VGND sg13g2_decap_8
XFILLER_28_372 VPWR VGND sg13g2_fill_1
XFILLER_16_578 VPWR VGND sg13g2_decap_8
XFILLER_12_773 VPWR VGND sg13g2_fill_2
XFILLER_15_1015 VPWR VGND sg13g2_decap_8
XFILLER_8_755 VPWR VGND sg13g2_fill_1
XFILLER_11_272 VPWR VGND sg13g2_fill_2
XFILLER_7_265 VPWR VGND sg13g2_decap_8
XFILLER_3_460 VPWR VGND sg13g2_fill_1
X_3260_ net1230 net999 _1703_ VPWR VGND sg13g2_nor2b_1
X_3191_ net1006 net1051 _1638_ VPWR VGND sg13g2_nor2b_1
XFILLER_39_615 VPWR VGND sg13g2_decap_8
Xfanout1250 net1253 net1250 VPWR VGND sg13g2_buf_8
Xfanout1272 ui_in[2] net1272 VPWR VGND sg13g2_buf_8
Xfanout1283 net1284 net1283 VPWR VGND sg13g2_buf_8
Xfanout1261 net1263 net1261 VPWR VGND sg13g2_buf_1
Xfanout1294 net1296 net1294 VPWR VGND sg13g2_buf_8
X_5901_ _1517_ VPWR _1518_ VGND _1513_ _1516_ sg13g2_o21ai_1
XFILLER_19_372 VPWR VGND sg13g2_fill_1
X_6145__129 VPWR VGND net129 sg13g2_tiehi
X_5832_ _1387_ _1457_ net1257 _1458_ VPWR VGND sg13g2_nand3_1
X_5763_ VPWR _0158_ _1392_ VGND sg13g2_inv_1
X_4714_ _0447_ VPWR _0448_ VGND net1305 net480 sg13g2_o21ai_1
X_5694_ VGND VPWR _1275_ _1334_ _1339_ net1251 sg13g2_a21oi_1
X_4645_ s0.data_out\[18\]\[6\] s0.data_out\[17\]\[6\] net1166 _0386_ VPWR VGND sg13g2_mux2_1
X_4576_ VGND VPWR _0323_ net498 net1302 sg13g2_or2_1
X_3527_ s0.data_out\[3\]\[0\] s0.data_out\[4\]\[0\] net987 _1944_ VPWR VGND sg13g2_mux2_1
X_3458_ net1314 VPWR _1880_ VGND net915 _1879_ sg13g2_o21ai_1
X_3389_ net994 _1703_ _1820_ VPWR VGND sg13g2_nor2_1
X_6177_ net94 VGND VPWR _0227_ s0.data_out\[3\]\[1\] clknet_leaf_5_clk sg13g2_dfrbpq_2
X_5128_ net1113 net1048 _0822_ VPWR VGND sg13g2_nor2b_1
X_5059_ net1129 VPWR _0762_ VGND net1228 net1114 sg13g2_o21ai_1
XFILLER_37_191 VPWR VGND sg13g2_decap_8
XFILLER_13_515 VPWR VGND sg13g2_fill_1
XFILLER_40_367 VPWR VGND sg13g2_fill_2
XFILLER_4_224 VPWR VGND sg13g2_fill_2
XFILLER_45_1019 VPWR VGND sg13g2_decap_8
XFILLER_1_942 VPWR VGND sg13g2_decap_8
X_6211__208 VPWR VGND net208 sg13g2_tiehi
XFILLER_0_452 VPWR VGND sg13g2_decap_8
XFILLER_49_968 VPWR VGND sg13g2_decap_8
XFILLER_48_478 VPWR VGND sg13g2_decap_8
Xhold71 _0006_ VPWR VGND net367 sg13g2_dlygate4sd3_1
Xhold82 s0.was_valid_out\[14\][0] VPWR VGND net378 sg13g2_dlygate4sd3_1
Xhold60 s0.data_out\[21\]\[6\] VPWR VGND net356 sg13g2_dlygate4sd3_1
Xhold93 _2534_ VPWR VGND net389 sg13g2_dlygate4sd3_1
XFILLER_29_681 VPWR VGND sg13g2_fill_2
XFILLER_44_640 VPWR VGND sg13g2_fill_1
XFILLER_17_876 VPWR VGND sg13g2_decap_4
XFILLER_16_386 VPWR VGND sg13g2_decap_8
XFILLER_32_868 VPWR VGND sg13g2_fill_2
XFILLER_6_31 VPWR VGND sg13g2_fill_2
X_4430_ _2753_ VPWR _2754_ VGND net1287 net410 sg13g2_o21ai_1
X_6005__280 VPWR VGND net280 sg13g2_tiehi
X_4361_ s0.data_out\[20\]\[2\] s0.data_out\[19\]\[2\] net1186 _2689_ VPWR VGND sg13g2_mux2_1
X_6100_ net178 VGND VPWR _0150_ s0.data_new_delayed\[6\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_3312_ VGND VPWR _1673_ _1747_ _1748_ net1004 sg13g2_a21oi_1
X_4292_ _2456_ VPWR _2630_ VGND net323 net1201 sg13g2_o21ai_1
X_3243_ s0.data_out\[7\]\[6\] s0.data_out\[6\]\[6\] net1010 _1688_ VPWR VGND sg13g2_mux2_1
X_6151__122 VPWR VGND net122 sg13g2_tiehi
X_6031_ net252 VGND VPWR _0081_ s0.data_out\[15\]\[6\] clknet_leaf_30_clk sg13g2_dfrbpq_2
XFILLER_39_423 VPWR VGND sg13g2_fill_2
XFILLER_6_1024 VPWR VGND sg13g2_decap_4
XFILLER_39_456 VPWR VGND sg13g2_fill_2
XFILLER_39_445 VPWR VGND sg13g2_fill_2
X_3174_ VGND VPWR _1564_ _1622_ _1623_ net1015 sg13g2_a21oi_1
XFILLER_13_0 VPWR VGND sg13g2_fill_2
Xfanout1091 net1092 net1091 VPWR VGND sg13g2_buf_2
Xfanout1080 net1081 net1080 VPWR VGND sg13g2_buf_8
XFILLER_48_990 VPWR VGND sg13g2_decap_8
XFILLER_25_18 VPWR VGND sg13g2_decap_8
X_5815_ s0.data_out\[9\]\[6\] s0.data_out\[8\]\[6\] net1033 _1441_ VPWR VGND sg13g2_mux2_1
XFILLER_23_835 VPWR VGND sg13g2_decap_8
X_5746_ net609 VPWR _1378_ VGND net1340 net451 sg13g2_o21ai_1
X_5677_ _1322_ _1321_ net1243 _1317_ net1237 VPWR VGND sg13g2_a22oi_1
X_4628_ s0.data_out\[18\]\[0\] s0.data_out\[17\]\[0\] net1163 _0369_ VPWR VGND sg13g2_mux2_1
X_4559_ net1169 VPWR _0308_ VGND _0306_ _0307_ sg13g2_o21ai_1
XFILLER_2_728 VPWR VGND sg13g2_decap_8
XFILLER_9_8 VPWR VGND sg13g2_decap_8
XFILLER_45_426 VPWR VGND sg13g2_decap_4
XFILLER_17_117 VPWR VGND sg13g2_decap_4
XFILLER_26_640 VPWR VGND sg13g2_decap_8
XFILLER_25_150 VPWR VGND sg13g2_fill_1
XFILLER_40_186 VPWR VGND sg13g2_decap_8
XFILLER_15_95 VPWR VGND sg13g2_fill_1
XFILLER_5_522 VPWR VGND sg13g2_decap_8
XFILLER_31_50 VPWR VGND sg13g2_decap_8
XFILLER_31_94 VPWR VGND sg13g2_fill_1
XFILLER_5_599 VPWR VGND sg13g2_decap_8
XFILLER_5_588 VPWR VGND sg13g2_decap_8
Xoutput4 net4 uo_out[2] VPWR VGND sg13g2_buf_1
XFILLER_0_260 VPWR VGND sg13g2_decap_8
XFILLER_49_765 VPWR VGND sg13g2_decap_8
XFILLER_16_150 VPWR VGND sg13g2_fill_1
X_3930_ net951 VPWR _2309_ VGND _2307_ _2308_ sg13g2_o21ai_1
XFILLER_44_481 VPWR VGND sg13g2_decap_4
X_3861_ s0.data_out\[2\]\[3\] s0.data_out\[1\]\[3\] net958 _2246_ VPWR VGND sg13g2_mux2_1
XFILLER_32_654 VPWR VGND sg13g2_fill_1
X_3792_ _2184_ net930 _2183_ VPWR VGND sg13g2_nand2_1
X_5600_ _1251_ VPWR _1252_ VGND net1341 net418 sg13g2_o21ai_1
X_5531_ VGND VPWR net1090 _1187_ _1188_ _1133_ sg13g2_a21oi_1
X_5462_ net1077 s0.data_out\[10\]\[0\] _1127_ VPWR VGND sg13g2_and2_1
X_4413_ net1183 VPWR _2739_ VGND net1226 net1170 sg13g2_o21ai_1
X_5393_ _1062_ net1099 net568 VPWR VGND sg13g2_nand2_1
X_4344_ VPWR _0020_ _2674_ VGND sg13g2_inv_1
XFILLER_28_1014 VPWR VGND sg13g2_decap_8
X_6014_ net270 VGND VPWR _0064_ s0.data_out\[16\]\[1\] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_4275_ _2614_ VPWR _2615_ VGND net1254 _2605_ sg13g2_o21ai_1
X_3226_ _1670_ net1005 _1624_ _1671_ VPWR VGND sg13g2_a21o_1
XFILLER_28_916 VPWR VGND sg13g2_decap_8
XFILLER_39_264 VPWR VGND sg13g2_fill_1
XFILLER_36_17 VPWR VGND sg13g2_decap_8
X_3157_ s0.data_out\[6\]\[2\] s0.data_out\[7\]\[2\] net1019 _1608_ VPWR VGND sg13g2_mux2_1
XFILLER_28_927 VPWR VGND sg13g2_fill_1
XFILLER_43_919 VPWR VGND sg13g2_decap_8
XFILLER_35_470 VPWR VGND sg13g2_decap_8
X_5729_ _1359_ _1362_ net1340 _1363_ VPWR VGND sg13g2_nand3_1
XFILLER_19_927 VPWR VGND sg13g2_decap_8
XFILLER_46_768 VPWR VGND sg13g2_decap_8
XFILLER_34_908 VPWR VGND sg13g2_fill_1
X_5968__48 VPWR VGND net48 sg13g2_tiehi
XFILLER_26_470 VPWR VGND sg13g2_fill_1
XFILLER_13_142 VPWR VGND sg13g2_decap_8
XFILLER_42_985 VPWR VGND sg13g2_decap_8
XFILLER_9_102 VPWR VGND sg13g2_fill_2
XFILLER_13_186 VPWR VGND sg13g2_fill_2
X_6002__283 VPWR VGND net283 sg13g2_tiehi
XFILLER_3_10 VPWR VGND sg13g2_decap_4
X_4060_ VGND VPWR net1294 _2422_ _0268_ _2420_ sg13g2_a21oi_1
XFILLER_49_562 VPWR VGND sg13g2_decap_8
XFILLER_3_1027 VPWR VGND sg13g2_fill_2
XFILLER_36_278 VPWR VGND sg13g2_fill_2
X_4962_ _0604_ VPWR _0672_ VGND net1142 _2486_ sg13g2_o21ai_1
X_4893_ _0610_ net1142 net554 VPWR VGND sg13g2_nand2_1
X_3913_ net940 net1073 _2294_ VPWR VGND sg13g2_nor2b_1
XFILLER_32_451 VPWR VGND sg13g2_decap_4
X_3844_ VGND VPWR _2230_ net553 net1298 sg13g2_or2_1
XFILLER_20_646 VPWR VGND sg13g2_fill_2
X_3775_ _2169_ VPWR _2170_ VGND net962 _2052_ sg13g2_o21ai_1
X_5514_ _1172_ VPWR _1173_ VGND _1168_ _1171_ sg13g2_o21ai_1
X_5445_ VGND VPWR _1114_ net1209 net302 sg13g2_or2_1
X_5376_ VPWR _0116_ net502 VGND sg13g2_inv_1
X_4327_ _2659_ VPWR _2660_ VGND _2655_ _2658_ sg13g2_o21ai_1
X_4258_ VGND VPWR net1204 _2597_ _2598_ _2561_ sg13g2_a21oi_1
X_3209_ _1654_ net1008 net537 VPWR VGND sg13g2_nand2_1
XFILLER_27_201 VPWR VGND sg13g2_decap_8
X_4189_ VPWR _0005_ net389 VGND sg13g2_inv_1
XFILLER_42_226 VPWR VGND sg13g2_fill_2
XFILLER_42_215 VPWR VGND sg13g2_decap_8
XFILLER_27_289 VPWR VGND sg13g2_fill_2
XFILLER_42_259 VPWR VGND sg13g2_decap_4
XFILLER_10_167 VPWR VGND sg13g2_fill_2
XFILLER_12_63 VPWR VGND sg13g2_fill_1
XFILLER_3_845 VPWR VGND sg13g2_decap_8
Xhold190 s0.data_out\[11\]\[3\] VPWR VGND net486 sg13g2_dlygate4sd3_1
XFILLER_19_746 VPWR VGND sg13g2_decap_8
XFILLER_18_245 VPWR VGND sg13g2_decap_4
XFILLER_30_911 VPWR VGND sg13g2_fill_1
XFILLER_41_292 VPWR VGND sg13g2_fill_2
XFILLER_30_988 VPWR VGND sg13g2_decap_8
X_3560_ _1973_ net914 _1972_ VPWR VGND sg13g2_nand2_1
X_3491_ VGND VPWR _1912_ _1906_ net1233 sg13g2_or2_1
XFILLER_6_683 VPWR VGND sg13g2_decap_8
X_5230_ VPWR _0102_ net508 VGND sg13g2_inv_1
X_5161_ _0854_ _0853_ net1242 _0849_ net1236 VPWR VGND sg13g2_a22oi_1
XFILLER_25_1006 VPWR VGND sg13g2_decap_8
X_4112_ _2471_ net983 VPWR VGND sg13g2_inv_2
X_5092_ _0790_ VPWR _0791_ VGND _0786_ _0789_ sg13g2_o21ai_1
X_4043_ VGND VPWR net1292 _2409_ _0264_ _2406_ sg13g2_a21oi_1
XFILLER_37_576 VPWR VGND sg13g2_fill_2
XFILLER_37_565 VPWR VGND sg13g2_fill_2
X_5994_ net292 VGND VPWR _0044_ s0.data_out\[18\]\[5\] clknet_leaf_3_clk sg13g2_dfrbpq_2
X_4945_ VPWR _0075_ _0657_ VGND sg13g2_inv_1
X_4876_ _0550_ VPWR _0593_ VGND net922 _0592_ sg13g2_o21ai_1
X_5955__62 VPWR VGND net62 sg13g2_tiehi
X_6083__196 VPWR VGND net196 sg13g2_tiehi
XFILLER_33_793 VPWR VGND sg13g2_fill_1
X_3827_ net962 VPWR _2215_ VGND _2213_ _2214_ sg13g2_o21ai_1
X_3758_ _2155_ _2154_ net1248 _2151_ net1255 VPWR VGND sg13g2_a22oi_1
XFILLER_3_108 VPWR VGND sg13g2_fill_1
X_3689_ _2090_ net932 _2089_ VPWR VGND sg13g2_nand2_1
X_5428_ _1096_ net1092 _1036_ _1097_ VPWR VGND sg13g2_a21o_1
X_5359_ net614 VPWR _1033_ VGND net1334 net472 sg13g2_o21ai_1
XFILLER_48_808 VPWR VGND sg13g2_decap_8
XFILLER_0_859 VPWR VGND sg13g2_decap_8
XFILLER_28_565 VPWR VGND sg13g2_fill_2
XFILLER_31_708 VPWR VGND sg13g2_fill_1
XFILLER_30_207 VPWR VGND sg13g2_fill_1
XFILLER_8_904 VPWR VGND sg13g2_fill_2
XFILLER_8_915 VPWR VGND sg13g2_decap_8
XFILLER_12_999 VPWR VGND sg13g2_decap_8
X_6202__66 VPWR VGND net66 sg13g2_tiehi
XFILLER_7_447 VPWR VGND sg13g2_decap_8
XFILLER_3_675 VPWR VGND sg13g2_decap_4
XFILLER_38_307 VPWR VGND sg13g2_fill_1
XFILLER_19_532 VPWR VGND sg13g2_fill_1
XFILLER_47_885 VPWR VGND sg13g2_decap_8
XFILLER_34_568 VPWR VGND sg13g2_fill_2
XFILLER_34_579 VPWR VGND sg13g2_fill_1
XFILLER_9_31 VPWR VGND sg13g2_fill_2
X_4730_ _0461_ VPWR _0462_ VGND _0457_ _0460_ sg13g2_o21ai_1
XFILLER_30_730 VPWR VGND sg13g2_fill_2
X_4661_ _0401_ _0333_ net1255 _0402_ VPWR VGND sg13g2_a21o_1
X_3612_ s0.data_out\[4\]\[7\] s0.data_out\[3\]\[7\] net978 _2021_ VPWR VGND sg13g2_mux2_1
X_4592_ _0333_ _0336_ net1303 _0337_ VPWR VGND sg13g2_nand3_1
X_5952__65 VPWR VGND net65 sg13g2_tiehi
XFILLER_7_992 VPWR VGND sg13g2_decap_8
X_3543_ _1958_ net420 net987 VPWR VGND sg13g2_nand2b_1
XFILLER_43_0 VPWR VGND sg13g2_fill_2
X_3474_ VPWR VGND _1828_ net1282 _1894_ net1277 _1895_ _1891_ sg13g2_a221oi_1
X_6193_ net77 VGND VPWR _0243_ s0.data_out\[2\]\[5\] clknet_leaf_11_clk sg13g2_dfrbpq_2
X_5213_ _0900_ VPWR _0901_ VGND net1332 net471 sg13g2_o21ai_1
X_5144_ net1279 _0833_ _0837_ VPWR VGND sg13g2_nor2_1
XFILLER_38_841 VPWR VGND sg13g2_decap_4
X_5075_ _0772_ _0775_ net1321 _0776_ VPWR VGND sg13g2_nand3_1
X_4026_ VGND VPWR net363 _2465_ _2397_ net1225 sg13g2_a21oi_1
XFILLER_38_852 VPWR VGND sg13g2_fill_1
X_5977_ net38 VGND VPWR _0027_ s0.data_out\[19\]\[0\] clknet_leaf_36_clk sg13g2_dfrbpq_2
XFILLER_13_719 VPWR VGND sg13g2_decap_8
X_4928_ _0641_ _0642_ _0643_ VPWR VGND sg13g2_nor2_1
X_4859_ VGND VPWR _0496_ _0577_ _0578_ net1148 sg13g2_a21oi_1
XFILLER_20_262 VPWR VGND sg13g2_decap_4
XFILLER_20_273 VPWR VGND sg13g2_decap_8
Xclkbuf_3_0__f_clk clknet_0_clk clknet_3_0__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_20_295 VPWR VGND sg13g2_fill_1
XFILLER_0_656 VPWR VGND sg13g2_decap_8
XFILLER_48_605 VPWR VGND sg13g2_decap_8
XFILLER_18_40 VPWR VGND sg13g2_fill_1
XFILLER_44_822 VPWR VGND sg13g2_decap_8
XFILLER_16_524 VPWR VGND sg13g2_decap_4
XFILLER_43_343 VPWR VGND sg13g2_fill_1
XFILLER_43_321 VPWR VGND sg13g2_fill_2
XFILLER_44_899 VPWR VGND sg13g2_decap_8
XFILLER_12_763 VPWR VGND sg13g2_fill_1
XFILLER_12_796 VPWR VGND sg13g2_decap_8
XFILLER_7_244 VPWR VGND sg13g2_fill_1
X_6138__137 VPWR VGND net137 sg13g2_tiehi
XFILLER_4_984 VPWR VGND sg13g2_decap_8
XFILLER_3_450 VPWR VGND sg13g2_fill_1
X_3190_ VGND VPWR _1556_ _1636_ _1637_ net1015 sg13g2_a21oi_1
Xfanout1240 net1241 net1240 VPWR VGND sg13g2_buf_8
Xfanout1273 net1276 net1273 VPWR VGND sg13g2_buf_8
Xfanout1262 net1263 net1262 VPWR VGND sg13g2_buf_8
Xfanout1251 net1253 net1251 VPWR VGND sg13g2_buf_8
Xfanout1295 net1296 net1295 VPWR VGND sg13g2_buf_1
Xfanout1284 ui_in[0] net1284 VPWR VGND sg13g2_buf_8
XFILLER_47_682 VPWR VGND sg13g2_decap_8
X_5900_ VGND VPWR _1517_ net482 net1342 sg13g2_or2_1
XFILLER_35_866 VPWR VGND sg13g2_fill_2
XFILLER_19_395 VPWR VGND sg13g2_decap_8
X_5831_ _1457_ net343 _1456_ VPWR VGND sg13g2_nand2b_1
X_5762_ _1391_ VPWR _1392_ VGND net1342 net442 sg13g2_o21ai_1
X_4713_ _0443_ _0446_ net1305 _0447_ VPWR VGND sg13g2_nand3_1
XFILLER_30_560 VPWR VGND sg13g2_decap_4
XFILLER_30_582 VPWR VGND sg13g2_decap_8
X_5693_ net1266 _1311_ _1338_ VPWR VGND sg13g2_nor2_1
X_4644_ _0385_ net1165 net572 VPWR VGND sg13g2_nand2_1
X_6080__199 VPWR VGND net199 sg13g2_tiehi
X_4575_ net1301 VPWR _0322_ VGND net925 _0321_ sg13g2_o21ai_1
X_3526_ net1219 _1937_ _0213_ VPWR VGND sg13g2_nor2_1
X_3457_ VGND VPWR net984 net535 _1879_ _1878_ sg13g2_a21oi_1
X_3388_ _1817_ _1818_ _1819_ VPWR VGND sg13g2_nor2_1
X_6176_ net95 VGND VPWR _0226_ s0.data_out\[3\]\[0\] clknet_leaf_6_clk sg13g2_dfrbpq_2
X_5127_ VGND VPWR _0729_ _0820_ _0821_ net1128 sg13g2_a21oi_1
XFILLER_29_126 VPWR VGND sg13g2_decap_8
X_5058_ net1321 net303 _0084_ VPWR VGND sg13g2_and2_1
XFILLER_44_118 VPWR VGND sg13g2_decap_8
X_4009_ _2320_ VPWR _2382_ VGND net928 _2381_ sg13g2_o21ai_1
XFILLER_37_170 VPWR VGND sg13g2_decap_8
XFILLER_25_332 VPWR VGND sg13g2_decap_8
XFILLER_40_302 VPWR VGND sg13g2_decap_4
XFILLER_26_899 VPWR VGND sg13g2_fill_2
XFILLER_41_847 VPWR VGND sg13g2_fill_1
XFILLER_41_836 VPWR VGND sg13g2_decap_8
XFILLER_9_509 VPWR VGND sg13g2_decap_8
XFILLER_21_582 VPWR VGND sg13g2_decap_4
XFILLER_5_715 VPWR VGND sg13g2_decap_8
XFILLER_1_921 VPWR VGND sg13g2_decap_8
XFILLER_0_431 VPWR VGND sg13g2_decap_8
XFILLER_49_947 VPWR VGND sg13g2_decap_8
XFILLER_1_998 VPWR VGND sg13g2_decap_8
Xhold50 s0.was_valid_out\[13\][0] VPWR VGND net346 sg13g2_dlygate4sd3_1
XFILLER_48_457 VPWR VGND sg13g2_decap_8
Xhold72 s0.data_out\[21\]\[0\] VPWR VGND net368 sg13g2_dlygate4sd3_1
Xhold61 _0009_ VPWR VGND net357 sg13g2_dlygate4sd3_1
Xhold83 s0.was_valid_out\[10\][0] VPWR VGND net379 sg13g2_dlygate4sd3_1
XFILLER_17_822 VPWR VGND sg13g2_fill_2
Xhold94 s0.data_out\[8\]\[0\] VPWR VGND net390 sg13g2_dlygate4sd3_1
XFILLER_45_93 VPWR VGND sg13g2_fill_1
XFILLER_31_302 VPWR VGND sg13g2_fill_1
XFILLER_31_313 VPWR VGND sg13g2_fill_2
X_6144__130 VPWR VGND net130 sg13g2_tiehi
XFILLER_40_880 VPWR VGND sg13g2_fill_2
XFILLER_6_43 VPWR VGND sg13g2_fill_1
X_4360_ VPWR _0022_ net524 VGND sg13g2_inv_1
X_3311_ _1747_ net352 net1009 VPWR VGND sg13g2_nand2b_1
X_4291_ net1182 _2623_ _2629_ VPWR VGND sg13g2_nor2_1
X_3242_ _1687_ net1009 net557 VPWR VGND sg13g2_nand2_1
XFILLER_6_1003 VPWR VGND sg13g2_decap_8
X_6030_ net253 VGND VPWR _0080_ s0.data_out\[15\]\[5\] clknet_leaf_23_clk sg13g2_dfrbpq_2
X_3173_ _1622_ net423 net1019 VPWR VGND sg13g2_nand2b_1
Xfanout1092 net1094 net1092 VPWR VGND sg13g2_buf_2
Xfanout1070 net1072 net1070 VPWR VGND sg13g2_buf_8
Xfanout1081 net1083 net1081 VPWR VGND sg13g2_buf_8
XFILLER_19_181 VPWR VGND sg13g2_fill_2
XFILLER_23_814 VPWR VGND sg13g2_fill_2
XFILLER_34_151 VPWR VGND sg13g2_decap_4
X_5814_ _1440_ net1032 net587 VPWR VGND sg13g2_nand2_1
XFILLER_35_696 VPWR VGND sg13g2_decap_4
X_5745_ _1373_ _1376_ net1340 _1377_ VPWR VGND sg13g2_nand3_1
X_5676_ VGND VPWR net1083 _1320_ _1321_ _1282_ sg13g2_a21oi_1
X_4627_ VGND VPWR net1169 _0367_ _0368_ _0312_ sg13g2_a21oi_1
X_4558_ net1155 net1076 _0307_ VPWR VGND sg13g2_nor2b_1
XFILLER_2_707 VPWR VGND sg13g2_decap_8
X_3509_ _1914_ _1929_ _1930_ VPWR VGND sg13g2_nor2b_1
X_4489_ _2804_ VPWR _2805_ VGND net1174 _2483_ sg13g2_o21ai_1
X_6159_ net114 VGND VPWR _0209_ s0.data_out\[5\]\[7\] clknet_leaf_12_clk sg13g2_dfrbpq_2
Xclkbuf_leaf_37_clk clknet_3_0__leaf_clk clknet_leaf_37_clk VPWR VGND sg13g2_buf_8
XFILLER_14_836 VPWR VGND sg13g2_fill_1
X_6128__147 VPWR VGND net147 sg13g2_tiehi
XFILLER_25_184 VPWR VGND sg13g2_fill_1
XFILLER_40_121 VPWR VGND sg13g2_decap_8
XFILLER_22_880 VPWR VGND sg13g2_fill_2
XFILLER_5_556 VPWR VGND sg13g2_decap_8
XFILLER_31_84 VPWR VGND sg13g2_fill_1
Xoutput5 net5 uo_out[3] VPWR VGND sg13g2_buf_1
XFILLER_1_795 VPWR VGND sg13g2_decap_8
XFILLER_49_744 VPWR VGND sg13g2_decap_8
XFILLER_36_449 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_28_clk clknet_3_5__leaf_clk clknet_leaf_28_clk VPWR VGND sg13g2_buf_8
X_3860_ _2245_ net955 net513 VPWR VGND sg13g2_nand2_1
XFILLER_20_839 VPWR VGND sg13g2_decap_8
X_3791_ s0.data_out\[1\]\[1\] s0.data_out\[2\]\[1\] net965 _2183_ VPWR VGND sg13g2_mux2_1
X_5530_ _1186_ net1077 _1134_ _1187_ VPWR VGND sg13g2_a21o_1
XFILLER_8_361 VPWR VGND sg13g2_decap_4
X_5461_ _1126_ net939 _1125_ VPWR VGND sg13g2_nand2_1
X_4412_ net1295 net297 _0024_ VPWR VGND sg13g2_and2_1
X_5392_ VPWR _0118_ _1061_ VGND sg13g2_inv_1
X_4343_ _2673_ VPWR _2674_ VGND net1285 net395 sg13g2_o21ai_1
X_4274_ _2612_ _2613_ _2614_ VPWR VGND sg13g2_nor2_1
X_3225_ s0.data_out\[7\]\[4\] s0.data_out\[6\]\[4\] net1009 _1670_ VPWR VGND sg13g2_mux2_1
X_6013_ net271 VGND VPWR _0063_ s0.data_out\[16\]\[0\] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_3156_ VPWR _0179_ _1607_ VGND sg13g2_inv_1
XFILLER_27_416 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_19_clk clknet_3_7__leaf_clk clknet_leaf_19_clk VPWR VGND sg13g2_buf_8
XFILLER_42_408 VPWR VGND sg13g2_fill_1
X_5977__38 VPWR VGND net38 sg13g2_tiehi
XFILLER_36_994 VPWR VGND sg13g2_decap_8
XFILLER_22_143 VPWR VGND sg13g2_decap_8
XFILLER_22_154 VPWR VGND sg13g2_fill_2
XFILLER_22_198 VPWR VGND sg13g2_decap_4
X_5728_ net1035 VPWR _1362_ VGND _1360_ _1361_ sg13g2_o21ai_1
X_3989_ _2362_ s0.data_out\[1\]\[3\] net946 VPWR VGND sg13g2_nand2b_1
X_5659_ VGND VPWR net1035 _1303_ _1304_ _1242_ sg13g2_a21oi_1
XFILLER_46_747 VPWR VGND sg13g2_decap_8
XFILLER_45_213 VPWR VGND sg13g2_decap_8
XFILLER_33_408 VPWR VGND sg13g2_fill_1
XFILLER_42_964 VPWR VGND sg13g2_decap_8
XFILLER_9_136 VPWR VGND sg13g2_decap_8
X_6141__133 VPWR VGND net133 sg13g2_tiehi
XFILLER_47_7 VPWR VGND sg13g2_decap_8
XFILLER_6_898 VPWR VGND sg13g2_decap_8
XFILLER_3_55 VPWR VGND sg13g2_decap_4
XFILLER_49_541 VPWR VGND sg13g2_decap_8
XFILLER_1_592 VPWR VGND sg13g2_decap_8
XFILLER_37_725 VPWR VGND sg13g2_fill_2
XFILLER_3_1006 VPWR VGND sg13g2_decap_8
XFILLER_3_99 VPWR VGND sg13g2_fill_2
XFILLER_37_747 VPWR VGND sg13g2_fill_1
X_4961_ VPWR _0077_ _0671_ VGND sg13g2_inv_1
XFILLER_18_994 VPWR VGND sg13g2_decap_8
XFILLER_33_920 VPWR VGND sg13g2_fill_2
X_4892_ _0608_ VPWR _0609_ VGND net1213 _0593_ sg13g2_o21ai_1
X_3912_ net941 s0.data_out\[0\]\[0\] _2293_ VPWR VGND sg13g2_and2_1
X_3843_ net1298 VPWR _2229_ VGND _2458_ _2228_ sg13g2_o21ai_1
XFILLER_33_997 VPWR VGND sg13g2_decap_8
X_3774_ VPWR _2169_ _2168_ VGND sg13g2_inv_1
X_5513_ VGND VPWR _1172_ net527 net1345 sg13g2_or2_1
Xclkbuf_leaf_8_clk clknet_3_2__leaf_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
X_5444_ _1000_ _1111_ _1112_ _1113_ VPWR VGND sg13g2_nor3_1
X_5375_ _1046_ VPWR _1047_ VGND _1042_ _1045_ sg13g2_o21ai_1
X_4326_ VGND VPWR _2659_ net560 net1286 sg13g2_or2_1
XFILLER_47_28 VPWR VGND sg13g2_fill_2
X_4257_ _2596_ net1195 _2557_ _2597_ VPWR VGND sg13g2_a21o_1
X_4188_ _2533_ VPWR _2534_ VGND net1285 net388 sg13g2_o21ai_1
X_3208_ _1609_ VPWR _1653_ VGND net917 _1652_ sg13g2_o21ai_1
X_3139_ VGND VPWR _2444_ _1592_ _0176_ _1593_ sg13g2_a21oi_1
XFILLER_42_205 VPWR VGND sg13g2_fill_1
XFILLER_24_986 VPWR VGND sg13g2_decap_8
XFILLER_7_618 VPWR VGND sg13g2_decap_8
XFILLER_12_75 VPWR VGND sg13g2_fill_2
XFILLER_3_824 VPWR VGND sg13g2_decap_8
Xhold180 s0.data_out\[16\]\[1\] VPWR VGND net476 sg13g2_dlygate4sd3_1
Xhold191 s0.data_out\[8\]\[2\] VPWR VGND net487 sg13g2_dlygate4sd3_1
XFILLER_42_783 VPWR VGND sg13g2_decap_8
XFILLER_42_772 VPWR VGND sg13g2_fill_1
X_5964__52 VPWR VGND net52 sg13g2_tiehi
X_3490_ _1911_ _1910_ net1240 _1906_ net1233 VPWR VGND sg13g2_a22oi_1
XFILLER_6_673 VPWR VGND sg13g2_decap_4
XFILLER_5_172 VPWR VGND sg13g2_decap_8
XFILLER_5_161 VPWR VGND sg13g2_decap_4
X_5160_ VGND VPWR net1128 _0852_ _0853_ _0814_ sg13g2_a21oi_1
X_4111_ VPWR _2470_ net994 VGND sg13g2_inv_1
X_5091_ VGND VPWR _0790_ net573 net1333 sg13g2_or2_1
XFILLER_37_500 VPWR VGND sg13g2_decap_8
X_4042_ VPWR _2409_ _2408_ VGND sg13g2_inv_1
XFILLER_37_533 VPWR VGND sg13g2_decap_4
X_5993_ net293 VGND VPWR _0043_ s0.data_out\[18\]\[4\] clknet_leaf_4_clk sg13g2_dfrbpq_2
XFILLER_40_709 VPWR VGND sg13g2_fill_2
X_4944_ _0656_ VPWR _0657_ VGND net1318 net461 sg13g2_o21ai_1
XFILLER_33_750 VPWR VGND sg13g2_fill_2
X_4875_ VGND VPWR net1134 _0591_ _0592_ _0552_ sg13g2_a21oi_1
XFILLER_21_934 VPWR VGND sg13g2_fill_2
X_3826_ net953 net1053 _2214_ VPWR VGND sg13g2_nor2b_1
XFILLER_20_444 VPWR VGND sg13g2_decap_8
X_3757_ VGND VPWR net973 _2153_ _2154_ _2097_ sg13g2_a21oi_1
X_3688_ s0.data_out\[2\]\[4\] s0.data_out\[3\]\[4\] net976 _2089_ VPWR VGND sg13g2_mux2_1
X_5427_ s0.data_out\[12\]\[4\] s0.data_out\[11\]\[4\] net1098 _1096_ VPWR VGND sg13g2_mux2_1
XFILLER_0_838 VPWR VGND sg13g2_decap_8
X_5358_ _1028_ _1031_ net1334 _1032_ VPWR VGND sg13g2_nand3_1
X_4309_ net1193 VPWR _2644_ VGND _2642_ _2643_ sg13g2_o21ai_1
X_5289_ s0.data_out\[13\]\[6\] s0.data_out\[12\]\[6\] net1111 _0970_ VPWR VGND sg13g2_mux2_1
XFILLER_43_525 VPWR VGND sg13g2_decap_8
XFILLER_15_227 VPWR VGND sg13g2_fill_1
XFILLER_12_978 VPWR VGND sg13g2_decap_8
XFILLER_23_41 VPWR VGND sg13g2_fill_2
XFILLER_23_52 VPWR VGND sg13g2_fill_1
XFILLER_23_63 VPWR VGND sg13g2_decap_4
XFILLER_48_1018 VPWR VGND sg13g2_decap_8
XFILLER_2_164 VPWR VGND sg13g2_decap_4
XFILLER_47_864 VPWR VGND sg13g2_decap_8
XFILLER_46_374 VPWR VGND sg13g2_decap_4
XFILLER_0_56 VPWR VGND sg13g2_decap_4
XFILLER_9_43 VPWR VGND sg13g2_decap_8
X_4660_ _0401_ net1171 _0400_ VPWR VGND sg13g2_nand2b_1
XFILLER_30_775 VPWR VGND sg13g2_decap_4
X_3611_ _2020_ net977 net515 VPWR VGND sg13g2_nand2_1
XFILLER_7_971 VPWR VGND sg13g2_decap_8
X_4591_ net1171 VPWR _0336_ VGND _0334_ _0335_ sg13g2_o21ai_1
X_3542_ VPWR _0215_ _1957_ VGND sg13g2_inv_1
X_3473_ _1894_ net990 _1893_ VPWR VGND sg13g2_nand2b_1
X_6192_ net78 VGND VPWR _0242_ s0.data_out\[2\]\[4\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_5212_ _0896_ _0899_ net1332 _0900_ VPWR VGND sg13g2_nand3_1
XFILLER_36_0 VPWR VGND sg13g2_decap_8
X_5143_ _0836_ net1127 _0835_ VPWR VGND sg13g2_nand2b_1
XFILLER_28_19 VPWR VGND sg13g2_fill_2
X_5074_ net1127 VPWR _0775_ VGND _0773_ _0774_ sg13g2_o21ai_1
X_4025_ net1289 net305 _0259_ VPWR VGND sg13g2_and2_1
XFILLER_38_897 VPWR VGND sg13g2_fill_2
X_5976_ net39 VGND VPWR _0026_ s0.valid_out\[19\][0] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_25_569 VPWR VGND sg13g2_fill_2
X_4927_ net1228 net1130 _0642_ VPWR VGND sg13g2_nor2b_1
X_4858_ _0577_ s0.data_out\[15\]\[6\] net1153 VPWR VGND sg13g2_nand2b_1
X_3809_ net950 s0.data_out\[1\]\[3\] _2199_ VPWR VGND sg13g2_and2_1
X_4789_ _0515_ VPWR _0518_ VGND net1262 _0493_ sg13g2_o21ai_1
XFILLER_0_635 VPWR VGND sg13g2_decap_8
XFILLER_47_149 VPWR VGND sg13g2_decap_4
XFILLER_44_801 VPWR VGND sg13g2_decap_8
XFILLER_16_536 VPWR VGND sg13g2_fill_2
XFILLER_44_878 VPWR VGND sg13g2_decap_8
XFILLER_24_591 VPWR VGND sg13g2_decap_8
XFILLER_31_528 VPWR VGND sg13g2_fill_2
XFILLER_8_746 VPWR VGND sg13g2_decap_8
XFILLER_11_252 VPWR VGND sg13g2_decap_8
XFILLER_11_274 VPWR VGND sg13g2_fill_1
XFILLER_8_779 VPWR VGND sg13g2_fill_2
XFILLER_4_963 VPWR VGND sg13g2_decap_8
Xfanout1241 net1245 net1241 VPWR VGND sg13g2_buf_8
Xfanout1230 uio_in[0] net1230 VPWR VGND sg13g2_buf_8
Xfanout1252 net1253 net1252 VPWR VGND sg13g2_buf_8
Xfanout1274 net1276 net1274 VPWR VGND sg13g2_buf_1
Xfanout1263 ui_in[3] net1263 VPWR VGND sg13g2_buf_8
Xfanout1296 net1300 net1296 VPWR VGND sg13g2_buf_8
Xfanout1285 net1291 net1285 VPWR VGND sg13g2_buf_8
XFILLER_47_661 VPWR VGND sg13g2_decap_8
XFILLER_19_352 VPWR VGND sg13g2_decap_8
XFILLER_34_322 VPWR VGND sg13g2_fill_1
X_5830_ VGND VPWR net1027 _1455_ _1456_ _1389_ sg13g2_a21oi_1
XFILLER_35_889 VPWR VGND sg13g2_decap_8
X_5761_ _1387_ _1390_ net1343 _1391_ VPWR VGND sg13g2_nand3_1
XFILLER_22_528 VPWR VGND sg13g2_decap_4
XFILLER_34_388 VPWR VGND sg13g2_fill_2
X_4712_ net1160 VPWR _0446_ VGND _0444_ _0445_ sg13g2_o21ai_1
X_5692_ VGND VPWR _1268_ _1330_ _1337_ net1257 sg13g2_a21oi_1
X_4643_ VGND VPWR net1171 _0383_ _0384_ _0354_ sg13g2_a21oi_1
X_4574_ VGND VPWR net1155 s0.data_out\[17\]\[2\] _0321_ _0320_ sg13g2_a21oi_1
X_3525_ _1938_ _1943_ _0212_ VPWR VGND sg13g2_nor2_1
X_3456_ net984 net1046 _1878_ VPWR VGND sg13g2_nor2b_1
X_3387_ net1226 net989 _1818_ VPWR VGND sg13g2_nor2b_1
X_6175_ net96 VGND VPWR _0225_ s0.valid_out\[3\][0] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5126_ _0820_ s0.data_out\[13\]\[7\] net1131 VPWR VGND sg13g2_nand2b_1
X_5057_ VGND VPWR _0756_ _0760_ _0083_ _0761_ sg13g2_a21oi_1
X_4008_ VGND VPWR net943 _2380_ _2381_ _2322_ sg13g2_a21oi_1
XFILLER_41_815 VPWR VGND sg13g2_decap_8
XFILLER_38_1028 VPWR VGND sg13g2_fill_1
XFILLER_38_1017 VPWR VGND sg13g2_decap_8
XFILLER_25_355 VPWR VGND sg13g2_decap_8
XFILLER_25_366 VPWR VGND sg13g2_fill_1
XFILLER_26_878 VPWR VGND sg13g2_decap_8
XFILLER_13_539 VPWR VGND sg13g2_fill_1
X_5959_ net58 VGND VPWR net357 s0.data_out\[21\]\[6\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_20_42 VPWR VGND sg13g2_fill_2
XFILLER_4_259 VPWR VGND sg13g2_decap_4
XFILLER_1_900 VPWR VGND sg13g2_decap_8
XFILLER_0_410 VPWR VGND sg13g2_decap_8
XFILLER_20_97 VPWR VGND sg13g2_decap_4
XFILLER_49_926 VPWR VGND sg13g2_decap_8
XFILLER_1_977 VPWR VGND sg13g2_decap_8
XFILLER_48_436 VPWR VGND sg13g2_decap_8
Xhold40 s0.shift_out\[15\][0] VPWR VGND net336 sg13g2_dlygate4sd3_1
Xhold73 _0003_ VPWR VGND net369 sg13g2_dlygate4sd3_1
Xhold51 _0097_ VPWR VGND net347 sg13g2_dlygate4sd3_1
Xhold62 s0.shift_out\[10\][0] VPWR VGND net358 sg13g2_dlygate4sd3_1
Xhold95 s0.data_out\[7\]\[0\] VPWR VGND net391 sg13g2_dlygate4sd3_1
XFILLER_29_650 VPWR VGND sg13g2_fill_1
XFILLER_29_661 VPWR VGND sg13g2_fill_1
XFILLER_29_683 VPWR VGND sg13g2_fill_1
Xhold84 _0133_ VPWR VGND net380 sg13g2_dlygate4sd3_1
XFILLER_44_631 VPWR VGND sg13g2_decap_8
XFILLER_17_856 VPWR VGND sg13g2_fill_2
XFILLER_45_50 VPWR VGND sg13g2_decap_8
XFILLER_44_675 VPWR VGND sg13g2_fill_2
XFILLER_43_130 VPWR VGND sg13g2_decap_4
XFILLER_43_185 VPWR VGND sg13g2_fill_1
XFILLER_31_325 VPWR VGND sg13g2_decap_8
XFILLER_32_826 VPWR VGND sg13g2_decap_8
XFILLER_32_837 VPWR VGND sg13g2_fill_1
XFILLER_31_336 VPWR VGND sg13g2_fill_1
XFILLER_31_347 VPWR VGND sg13g2_fill_1
XFILLER_40_870 VPWR VGND sg13g2_decap_4
XFILLER_12_583 VPWR VGND sg13g2_decap_8
XFILLER_8_565 VPWR VGND sg13g2_fill_2
XFILLER_6_33 VPWR VGND sg13g2_fill_1
X_3310_ VPWR _0194_ _1746_ VGND sg13g2_inv_1
XFILLER_3_281 VPWR VGND sg13g2_fill_1
X_4290_ VGND VPWR _2628_ _2627_ _2625_ sg13g2_or2_1
X_3241_ VGND VPWR net1018 _1685_ _1686_ _1644_ sg13g2_a21oi_1
XFILLER_39_425 VPWR VGND sg13g2_fill_1
X_3172_ VPWR _0181_ _1621_ VGND sg13g2_inv_1
Xfanout1060 net602 net1060 VPWR VGND sg13g2_buf_8
Xfanout1071 net1072 net1071 VPWR VGND sg13g2_buf_1
Xfanout1082 net1083 net1082 VPWR VGND sg13g2_buf_8
X_5989__25 VPWR VGND net25 sg13g2_tiehi
Xfanout1093 net1094 net1093 VPWR VGND sg13g2_buf_8
X_5813_ VGND VPWR net1038 _1438_ _1439_ _1408_ sg13g2_a21oi_1
XFILLER_22_303 VPWR VGND sg13g2_decap_8
X_5744_ net1036 VPWR _1376_ VGND _1374_ _1375_ sg13g2_o21ai_1
X_5675_ _1319_ net1039 _1283_ _1320_ VPWR VGND sg13g2_a21o_1
XFILLER_30_391 VPWR VGND sg13g2_fill_1
X_4626_ _0366_ net1156 _0313_ _0367_ VPWR VGND sg13g2_a21o_1
X_4557_ net1155 s0.data_out\[17\]\[0\] _0306_ VPWR VGND sg13g2_and2_1
X_3508_ _1922_ VPWR _1929_ VGND _1924_ _1925_ sg13g2_o21ai_1
X_4488_ _2804_ net1174 net498 VPWR VGND sg13g2_nand2_1
X_3439_ _1863_ net915 _1862_ VPWR VGND sg13g2_nand2_1
X_6158_ net115 VGND VPWR _0208_ s0.data_out\[5\]\[6\] clknet_leaf_13_clk sg13g2_dfrbpq_2
X_5109_ VPWR _0091_ _0805_ VGND sg13g2_inv_1
XFILLER_46_929 VPWR VGND sg13g2_decap_8
X_6089_ net189 VGND VPWR _0139_ s0.data_out\[10\]\[4\] clknet_leaf_21_clk sg13g2_dfrbpq_2
XFILLER_41_656 VPWR VGND sg13g2_decap_8
XFILLER_13_336 VPWR VGND sg13g2_decap_8
XFILLER_13_347 VPWR VGND sg13g2_decap_8
XFILLER_15_42 VPWR VGND sg13g2_fill_1
XFILLER_22_892 VPWR VGND sg13g2_fill_2
Xoutput6 net6 uo_out[4] VPWR VGND sg13g2_buf_1
XFILLER_49_723 VPWR VGND sg13g2_decap_8
XFILLER_1_774 VPWR VGND sg13g2_decap_8
XFILLER_36_428 VPWR VGND sg13g2_decap_8
XFILLER_17_642 VPWR VGND sg13g2_decap_8
XFILLER_45_984 VPWR VGND sg13g2_decap_8
XFILLER_31_100 VPWR VGND sg13g2_fill_2
XFILLER_13_881 VPWR VGND sg13g2_decap_4
X_3790_ VPWR _0238_ net425 VGND sg13g2_inv_1
XFILLER_9_874 VPWR VGND sg13g2_fill_1
X_5460_ s0.data_out\[10\]\[0\] s0.data_out\[11\]\[0\] net1096 _1125_ VPWR VGND sg13g2_mux2_1
XFILLER_8_384 VPWR VGND sg13g2_decap_8
X_4411_ VGND VPWR _2736_ _2737_ _0023_ _2738_ sg13g2_a21oi_1
X_5391_ _1060_ VPWR _1061_ VGND _1056_ _1059_ sg13g2_o21ai_1
X_4342_ _2669_ _2672_ net1289 _2673_ VPWR VGND sg13g2_nand3_1
X_4273_ net1246 _2609_ _2613_ VPWR VGND sg13g2_nor2_1
X_6012_ net272 VGND VPWR _0062_ s0.valid_out\[16\][0] clknet_leaf_33_clk sg13g2_dfrbpq_1
X_3224_ _1668_ VPWR _1669_ VGND net1212 _1653_ sg13g2_o21ai_1
.ends

